`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Eu/u28xpTcwH9/vC6LyUXt8zh+G6Z1US5rEInaWFwJ68VL9D0JZA+rGS21luLiZ9fpl+gxuCs995
+cZ4fAtijw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DgEZ3NGiCfrs93LCIy0I9taJ1U1Q7IJBxYKahP26GMUUP4ekQ/62YVqc/0mxvYPOT+3YJ/vLrSZM
Wk/OaPO0Y82IypIwxaqVMXsWCxsYuUvfr0TDfb0bbV4AnwY8GADD56ucrl1kVPlD/UmXpqzNXrdo
hCb2HZo5wizwAAtL9QA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LLu1gCxFf9Pk1NQMLzsAzeouO9NwyV88fRLhZMqDMdL3gj2EtZ47rLvU0egOr5WPncmgeACbVYtE
+Zhh3+YaWFu4rPV2URl/S5ZrwA1qca2nRHIMcnAkWjCftl96I51Hn4WNyYZIet9db+pXabZdq+yt
nQq9KPE9qwRVdsDliEpyv2Xzk5WinsSqUfBdTVjYqcFNsetruEbtGwR8tCRvsiFdKtsK4U6RvYQF
AQMgeSSwMaerguDAvJtWqnMtgh4wL8EhZbgB2SiHL+n7r32lOkVQ/I0i76qusMMt9yrNQ9y+/dWT
kb4gaMhXRYBEcrR0h8LSMIOA5MmjjXaTXLZ4nw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZNL0dpmy1SqdTTF+kaD+Y9ZMAshEOjbujfwUwmxTNJNu/MV9cdMzJH9uzT+3w6mydMsPy209HNuQ
1osPOmBWn8jlEBt0GEnAQFFyIC6S581InXu2c+Cf6jFs9NGR9zOsig8ZfPNV9js3dCnJdipW21DC
WtdTQZPmjPpClKufyG9ggZjoLI/y/lusVQ+PO4lxDfDhep5pUKErRA2+OTjRhqGgGqbl10Uf8Za+
oy1Wymwx2V8DvqnP9fCu645a5uywZQGuMfT86r09SVgzw5mEr36FVGCVZo8VtAKwReX3kfEB9y18
eATvhQw9qYOPxufoUF68SIOqRhdiXp4lva0Paw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mw3vH4Upj+FJlAT6nH2kJgBI26lJQHagQ7e4/GO2fLtksnbOWiqFSS1I+x1eOwgEwhUoviS22D+x
VtG5ece54r3oj/xJg9qOHoGNRjx/RIbZe7WP+4CO/ALn9DJn1TX6c2Xozt3oOwegD/GXTJNuWSSE
13Oy2h8+gqxBjjrDJso=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kcg8H/3QivWfQfyGC4SYEqxjl7e2cWjC0A1M8gGCLVpZgLscc9L3QEhQ6x9uDrpoPDv2agQTdxyD
GsltKDE1zrhjAlebTSMXpbP2+FAFg5vL/9a71PBxcfGIpdfFm3vNbdz5lE9ZpjQhHqV71REvaS1n
CCPuvRorvTH5mzDzykUrVzQFZ6qgs7QJotpFL1YdYU92uTKErW5gBUBA8aVQVySRnvVDV5yzeUeP
8IITfhhUSMI6ixPedUIT+Zi+cMh9t2rHZU8ZDTszq3isF7TeFlrjoJnxUmt753vj+YUJM4hcDRqa
ymYNwDX/kE9NQgYBaIcRzXuFGeu5zHEHHnERWQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LZCC7eP7l1dilV3mDVQO3ND+JpbIpGhQ6xrAhA6ocE7h9pcPJtXySWQFQYBiq7YMFy0utp1qPavP
9CLfYoD9inToGylGedB7CZNDAmyvtL5d0n8c0Aemql9BVkFTwFeVCaRPiBVEyPP40QTuZ9Sy0ia3
doTdkiGfiUECwTy8F2kOLR3rrHLWevI8WyiL8wQKX+3FBRT9alyCkwepi8B6TeI7XusjuGVKHLEU
/jiDTw7icrV9nbNY+q1Hqy6d375V3fYJlJVC96/bgh5q5pg/SAlylUE0zH0mD0FbuO0WSKR/4HEK
UBnGiGSayXwL7idxdhs74sbxk4BDPbiAbAxaiQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OUDR7dr4Lw9t82qyRv2xYFkNWwGByqtEVs6zx48AjeBh8DWa27osVoolvoyS3yHqzGPhgZS6idHk
4qQi3obLoyZPEE/bSGpI/Oo/FPk/DPpGr3KG5fZ+T5jtBRaDqncCZjv+GRx2MiuqsXi3ryP3Cx+e
wqEg/nhHi4/O2ITfIr8yixhji+WsLyRP9hKqNKLC5Kvl2A6rXfAnTI7Wlf4PT5HXs/mDoiqUYcsM
NVvZyWHqo2AOvksJA0DRh4f1+fMHQkEN92uyNvIS2vhSDvUtzVk3/T9rZWpXCVXmhjQGsWSLlwck
UwNrIXiksowKFpzZKy3eGdxZ7PuEDOFeHYPSDw==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p01Je5W/grzMYn5GLpSLOEMPYy5Dms8MjvO7R6xg/Co/k6hM6q+1KREB/v+Uzsw7XzHAu8PNgSOo
Di5wupKBN3prB8HLLzTdw8/JM3396y9hlcodNdj/eRDop9efL6o2wZekw3IGUxE9iSSQg0AnksfV
b5HCgGjbKj4qz9jQBzqca68gz0naWvEf3nHjclQA6x0wPaEDBqbnzn1z4VSfGiBe1u1O+FhiKcqO
ot61ms5Azfj/IM/HRrRgerKyCXivwiaW73EhZoSSm7QXAW7xCWgogbqB84+avMJ+ES3JGTe3jIEI
0zaqOODhLf3Dr0CVc5aohvg4f04vpot2YBo9Tg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 681264)
`protect data_block
rY4ieL5jQ+duq7sz0RxtGtoclBmI2IClsWJugx0T7u3Q46CIJyYSaycPjpWlWvyiGvjzGZb5bI+7
pH62wR02SfCLTbi+mSUygctVFW0jEWHdpcjV1D2/+b2FP1rCaJIs1VuJ9U1eacYXBMDPViaPTAtL
TYYDz3E25Oj5yf6/qRUvhvzUDsnWElNbXCGdiIZ73LpRfQ7u7v3Xy5w4mh4x/icxhXhtOP3b5BhT
jn0AjfJRdHa0EI+XAQ8LTrhT60nnDh9y8Kwx82V1Or47/2eupxMwnUC/I8mQE/2yJGXaSXqEVnug
YsDJoUSKJHD96dyB2GtfLHepM9v+En1tBllohr3/WFQnADkA+nvtYlJFiwtquBE/TG5RuxFmOLOX
T0x5UAMu36DPYulTcj4/wbBKxdYqXEQy0SaecYuMZjW8/t5k1T2ygfH5umim54ZuWNVp7RbJOGDW
+sBC5FitcbkvG/BOnFVV0AKFDAi6h+cJbrFFJIpXh86FW1j3aiWCtESbNn9u3Xeymm1SdfKcLEPu
dkzQj7NaeRcgqzt1HYhYtJ+sXa8xu8Acnoa3skOZW1AJCd8wB0dNMw4Y3N5lySL9KCFuGHroNFSD
j8ygBOO1oYEHCbFDGhhs1hAEO+5cyqhvUYnmM6dqj2YEajtV+6eccsB+TYqykIl9A3EFkBE6v8An
+hQ75LV4eW+FXpwme5UmdN0o0mTP2vWXTcOVig7PFcgDmYrl0bUTsX3+yjni5oonfGdnloL1zZkK
pnwPKSijYDwYl2o2p18PH8w6jRq/vvgjOfN9+6zB9c9twIkFxpsk2gQcAlKIOpxgls2Ha6V0C3bF
34F5Jvtss3GftzWUuT8VzNpKRo+YpITbpJAY8ikpPWAjwrYDMZ6+1H+z3JyjWCFn9iSNtgd73JEX
rZiDZW4cXFhcFRPM2ZCoqcpIfIQXVTjXqPSRz9JM8o5kQuz3cRu+Qo8iXvJYTiYI0U9Nvv02C3fp
276TKr+fgoN//x5aEn+Ys1sOtaKzm55gdjThbAkH3+kaTBg92O6VFDLk8J2wjQJ3hOTdE7FnzmI6
6N6ON0/Myxa58lAYl9UPfA0Jb3uOS2tLyCcS6uGB1hRXXwn6L8y29udI6JghbHbsayJyDvcoR4Ko
1NgtPiNiLmIayCTaPHab1kp/ZZS+UqPZEdByTuuOCxOTHB3gsivUoLqpbC2rIaNbkLw93CKNgKJ6
+NyNW23ICAy5odWxdvSQ7h7dxlCYOcLt2oriom7XL3f6kZeJL4GaqGzGl04Gw6/JCYCEB8xDnElx
mkutvSvKfJHT2Xkl0hMyyR6nJFa++oDnzQrkjLJYWe2RHBlDWsXxRZclge6cA9TbU5roC5jvBOL8
RYinAG3/N0CPkQ/uSKwLTsOJiIl2HgaTVVLWGr2HvFuJF0MKzSAA7cdxTCBq9wewhOfjI3HWbm+n
Ysx3GYvmje1QiepVL8c/zuWCYX7zIeYadNFF5XailhsBGVobm6Xnw0C5+Hm7bBy1n1a2iD99uiKD
feeyw4QWVTz1VqrcEz2FsmJuHSaBDaYuPWXI4yTLDeGd0j81zEqPrGWN0VPUnpKMv10pgIua510i
7N9LpbRQxebjSUQtt9/IxNODmTw/v8jOQh7YOwmUFBowzm4de02xw+0SlqZ/4VHi7MpKzA0Bpcq8
xDAc70sVPtmOnaoeEUf1TR+TqGl6UaVdoMIjcT3U4uWHrDmLCGfG1ckp2RSIvd2XrEJekAMHLBY4
gXYdoc/so7HS6ShlBOLepeOTd6KamamnVXGIRH2+kAJrZNO7U4/YRhr7BeiZ94nqRJIN3IOgr675
VyPiDIit1YgoW/MpZzxMFbJLLNpy4Uip4VPzy+O5dbPCTupU6F7zwRR6TteMH4l1eOUThVpnqhBY
Pa2rMlpbZqPpjG6Da3Jp9TRi+Y/dq+EuiNKcW0HlSlOYIGv8v6dD+7O9QFrJZWJpQWCPURE2Ipwt
8jCh/3Qr07AfdEnVzDc72Od1Uh1uAOjmPCaBkTpCPvDDYz8JEPoDH3Cl5Ke/WOLn9XetRJ1ttJ3z
iigwSKsZVkuugZsymVeak5vvh/jAia+ME9w9p8y0faeQgKuksysgnFy38DsRW5+Lt7VuCuOHxDaZ
eeYKPgVJEBahp3jb/7VRWyAt0qsA2IxkPt93/RnXzsBG0hNXci9TVrbtBtqbT0ExG3CKdTyA6qN1
6SbfyomIFwT4WKn3N7TCjAY+ayRaC8KRH51dunIrMCVXFEdYYSJ4nk/W4f+0gKYL59vNCMQZ3tBO
PCu1DX4Ew1BLqnk5LLgtTSkDsg/yZltsg0TZFexfXseliOaGfF5xC/MuVyQn0LARfVGvKVK0mrz8
vfZG4CnI27htjy3Y6K14+rxE9pQt7svFbNZBLnmMrwUJQgdZ7nvQaxl/yzu1NJFsxVPB+wi7kRXc
6TRsok93T3QkqEcOAQOlg3JBRB3SlUiDOqfFRwUyrWEOrW6HRZQz4jNuHFympUrZDKEuPRI1oMdp
2q1yTwYn4bQzfKfLbz5XqVQLB0hXgOJfnjP9sT+QnM/N/IT8O5Mr6abAlD4ijOAM0Z0zdUDDcGpX
JlSqJgnHQ8FmTFqDO6a/1fda2e+RPfVG0NTH3WEXc1t0QvPiiKynUG8Ev2Qu23Q84HHwzfuLkhRU
35Eh/BFTNKxdoyTl7iuL5xl5HKEumIhNFdFch13fckWplkqMHKnhk4WApDBmA0LOvqz191Cqa0D6
Y5DXaC1FxrHlMjQE11ED55Si8ro/rxK9sbiiPgD4F6plSVY6ZaywI2c7BnMEQ0M3B85ab/ubi4th
1qvabRdDSTFRb+vNhSJlkpEEIuFS5MAojy5bfn+bfS0l6RTs7p5b73XQty86zLBcc8qDj1RgQ01l
YXD8GUObDX0Jh4r1bVLF36Mvrn4ED5qbBnGnkc5ivlx5wY3CJCmWkn9edvPtFaZJ/9um7rJ4fZqa
e6ZXalvT+UiwS0r+pQ1yZzvlQRAKSamFZVU4uOmRfCiqAMvLogHeEMRQanPHtlRJt4/bywHUq5iC
r5t65hn9Q5c7izkyakSXwjDUG0JYhS9a4wJCmgvxrI18EQliPfnW7hn69/gv7b6Wu2BEzDU+2uFr
TaFNqNVhzB7sF/DD5DxxwzJkkG0d/dmw8SAjC7aM/lis/XIxKO2geOw7g3HxxbOBDviUyzDvmFW8
251j6t+Yka1phAg9NJA3/ls7/0v7Fk7z+2H+VULXA6tuSMkx9EloPi+gixR+h+wfqqvpDn902Bwh
tv6bJDc6dmY3U0yH9HA0E8Gk0a2kE1R/VG9rNmWFL3c8IJOo6AkH77FMdeZEM5MdMkus3O+iL9Cd
pRGUb+3Ia4qBBu6g1wd9ITUu4SzHgNndx5WlhdwtEw3B12tVQctu6hrz/zragJyG1oGMG3sC8oUu
TXhof1IABFZhwshVWn+cqwTgaDcQKZbyf2Q+nfoANwjeRvP1MoRaLkYV8+2FcPRwmlfUYyLq/rIX
tUYk0G6c0ag0179U3EN/l8DqGFRHAokYYtNXBC89DrazCCIqNUtkPnDuWbMw5rcNIbfSjB3UMx7/
wbW4wECfd/Y5LE6DIluaN3/uzqLA9GaCgcyqiAprzspWA/y32mVxFLWzVRqGhRn8u7mLaxbfk5ui
GxkT+drcSVLCneAiz6hugy73my9lSPHW7otTy40MB2HbZgk732Wjx/dowyY5ak0/FC8pfdH7huhL
2xeR9LEX3A18tLJtXrdRbMIkGBW5L6yXd1PocckXYGpHTEZPOPG9oD2KiTfa7NBK1mhKedZjxsCc
/YYr0bLbSHpzu5P6lUneWku06pIJIY7fVppU0K7gLsY0QsVlUdDSwWXRkSTZUSnQmfvTBBflYm2z
2pmwsWu904yCYFqE+Y6MzQGYT2h5iOTP6kBPbgbfHqDh2jqj+UdOgKwDr5s8VmXYj5bMpYoyhFPo
VZOJQvy4MTFPBz3YEPfnHxN+GQcPiUBfqNCtKwy5xYk65pNUeu5eoycV9KoN5cj6RQiYLcaSZl8O
uM7VGJbY3+EEXLXGJbnH2xOZoiuoAF4Xb85WqPYxcvKu5QmYE0FxL15PfahXw6wTLvKRF3fNLK2E
EF1yuRLrnOjlNGjVdpYt7FwFcILLqmlB+guCoLrfJDS782zXX7xxrDjA+qDktwEPmoUA84Vsfwh8
tM6yIhonOwVvdnCZYOKMA7w9WF5zsTKKgdPpuXN6U0S+reAW2/90kaWDZtM8zBjs4ct0Efb2P5eK
XvBPQE2ybf9QYLnSI2mMcT/wNLSdUzrVMBCU555HLa35sAdtqYLxGntdo6gQtpm58PhEJgNNPutO
5JHo8HQeDMhuf0H7IINN20A7MH8S0GPtERBW3l0dk+kzdVKlTa6Ht0rp9TH3Y/jQkpeVSJzW+C0p
i/WcoZopQOF0kbS6t0Eh6ydY8Y6OZHFZdXEQdSzVeBIuv9ARbkioL1O4k6xUp5Irau4Oq1OdDlQw
5hGaPVKOGPFoAwlGf69+4ExpFqKXjfPXDP7WcKAlxUpYuQG1Ewdp5c/040ujHTSvlpqVNBK5GYm5
cnz6jLGcSjWTh0jcMLhz1Upl6ngMp2P1sCxiL5gyf+/0YG5VELrTC+C5shUVPk12CC+iHfy6iDd/
k3sEyX515mn633dBcfwGyugZgvbnWIC0DCOpJX/QSwc2uW+Hf8KfJrQrU1/shIr61ENLXT9Jp3Vs
srrcazX1wR3MvnlQab/Cb+0RMKAfD9jToXvMI2TRyKrk8ieNiytLtlKjmpyxHz6JIl4dgTBDWddY
DoVBoOW0jybaBA6bdT3p6TJvf5QExPP5Sd42VzMXMw4/zKY8biIj/Si6nywp/Uq9eLqmJUVJysAJ
2lvrfu7ol/2QnwigwkUWZT1DbZYMkOB37B2ta0o2KmGINgJNdsIAVeX+xNf/J8AueKryCyKs1fe6
g8Rvo8WBX09acDJJI1f5HgQCY2SgKpISGhnaswewep/A7ETi54CA6ZvcUesYvGLw6QXNNlvVq7rr
z19vlh1CGEcR4ylGvmE1RiPy8C72jkjObyqv8+CJhDxeydZrZzUYAUWolnaeqf+7y6bgdjWR0Nlt
NaCk4bRTMk/ugqt3ypHcSbvaLFek/v8coHRFKAHAzCOKThX67owkQyA3OgJ7zwNJyKdBswDR+Kso
KFxDTBPta/AcLROI6q4NXRNQ7a8fav8HTR6pr2Z0PTb6QMz/1c+Fi5zyjTZdvIUQD9anZC7fm+gc
ET/5U3P3DbBdrQ+jF4IXeas8v4NhBGRHgGN1UmaXvg6Y0K9HbJcwBbw30hYaFjZHq1HTeo7E+Qka
zgzquvHsROtwyyP90NnqeHWxWCaj5l4UKjoqEQ1rL+LS45/t/V5bu4vfRJNsluhmmy/aveUv/9/s
kYukRVamGlecTq9fyyJAI496q1G+rTznytxIzcp334pPLPECSBLJ/MyVWq9a5a0j2Lmp+zCxMYfu
SDkrgzltVNOwuCYxAQxqlQIzN+s5iagTbLZpTsRVLvTVUQKz3LAaqd6JhlaQegc8pJrl+kS9OA5g
ZI9PZgUSReiqi7CAIjNz8fq1RP4y3IAU/e4i6BJXALNTBUkheZGNsTWwitz8SFMXCYMcZK15EwcM
+3MQYQ2mrcK62JS+O3HjwOVLFNHHOXVHLzh1eH5A7Gb0Okf+5S3Pi8qgpYckqQT6nnWhk/1oRROV
w/f6Je9LVZgAaV+UGchDz2a9cY0bRSDmpLiCKpulWIs3T10kuZRozicSevamBeV/acKRrStVFa1B
2KRSqQ0nKKgqxuDoKQ3ktRu9MdJpjk6ASJV8JyPFZPQfUtS6TyLt+sxkMavkj/Bw6gUB+38MUUbf
jzIM+7tQgRLjh6vkaggSsIpu8TwdVLRIgKsgBMZaIwbiuWGsyuSbVxJ/PSJjxY5q7rbfxI7ToIke
5MRIzpX+SqLPkFpKwMmcEkGXFcLm5d6AAQhLkWj9oftCY4S9gsNKPbzK+MHbpvXKRwTP6fRPTDtn
g0TM7jwI/YBBMxbS1dfvhvit//4qZZ4WVwNFmq2B7Qh2kOVUE/qvLg4ht/tthnjB3GuY2ELrRQnz
iHxOUCeMk1YeLZ8fQMzd6wA0U9P1R061MC6qXBW88tMcfizo9GPX3FAbz2Uu4bSXrrBC9G9SczXH
FDB8eGTKM15yCFMkzni0cfNWBd5jncpyrqcdwlOjZx2lUMnUGYxXHpcQlZdcWAumF99ru/LdJW4q
qVQPrDIm4+DpmEfA/6X9MMQWFMeYLjRPGEMbS5juFe2QGyI5TavGzAMkgawRCnqhTc6wvkwEPLBq
dKsvvIXUh7vg+akkMQ1Hi0hMbap5VZraHbPIaFp9IwxhYLIDIwpG+6MqwLwBJJLRG+33S5KBgS/x
HCm8hDq8yS/7wfeeNuDzFlrI35jEBukS3lZjoUWTsEEELttdramWyKIWWmleSfUp71uNHYU4zLrQ
dl5GEE7W0LP7zyUXV2WQhejY4Kqtf35bLPosiZ3tPLSjY+y4G7J6PiWMD1AWEtshHC6z+69Tq0Av
jvyeEs76KP+1zZ6oy3jI2JSOhQHLhifJerB40fDfXaiIgR0Ds/HCZFUyDglGBtbPhY9LQsCaKRtx
7MfoP6TQCGdbNqiJYAqPSfj+cErdIEGQJm/UEuFai0HSbONZSDhFDLz3CQhXdRHWGITpeDq8pcVo
X9JruCCtrxkr1S3qHa7V8LrrG9+oJfcNSvYF1fNAvah1DSfcXchtt2mHACap6IcMEwZukksPOpok
JL7X4ms+fueHeJSGC6CS2AeAtS8KWWQdUzmmcrIlgsbWxHDkCSbF6+2UTbGJSfojt8vuAfrUj42s
jAdZIEUnyj4RYdciNEOtSMZgQCAViEZsDJNnn6UMP0lyvXa/Ae2UL8U47wiFjoATtsjC2IieJ7vK
8jrFDgkcPbNrN+DzF1H+FodiNRYjTl9JZ5Ha4RKEYzCtA1bSD/FKeLy9GEFprwvaEauwpDMgkG3U
dvPFZ6Kdn7zLe9Li68CD1QKxTwICDrSVuLQ+jX7MGjgwx6d56k1NyN0lbjzSZWc0mmHCg1/M6lRd
Z7ZNCiIXctSQviqCpQh+cdn9+P3VhUzNUPcmEWUJ4C1yGJxVo62R+X0h5rUHF1GuRT1fSTwaSrnw
Pmy8Hl9cJ6969ugUiKOLtrH2f/IlxVwh92sBtNO/c11WcKgzlggkG+CDVwE3+n45iKt0P3jVSOqk
ilEiukQvny02pn4Ruj1R6CtjYl4UtTZX3tZFOaRWhPt33CMIaLt69Vw0mIc0dJbjFaXke1PjEAjD
LVgm3D97QyQNAKqu6swIbX9kN6s/j4OFQP+u7K0O1V78ND0KTm4xWMgbZavk+ThNvUeEJ2mh4g14
rP/ZTQz6rQZ5opD6sf2XBHtw7dx/OlONQqgGbrkcV/Z4Yp8BRw/UBZO4N1V2HZ0LYtjXI9dQaBXa
ysjTgKfZe9znAjGAZ83tygBWsE8z3EJnjiBXGL5XMBEv3o8c2DkUoblbksq/d4LnfSJF4T1ghNt7
MlHFQ4i9R8wK/at3IuOHMdgFPBoBfFY7igLNjghOF0bBH9KjleA8/CX2QAnAmY8rB1hYg/7O9aQq
wxMNQEwA/bOm/wpBye0TRJ/1tvym6h7kzFe6FbpbIldoIHqLrwG8jpcYXnaTT+F1PQ/dd9kYIoLl
TrIcMv9QMMSpQyqU5S8gB4DKVXXWxnvjLvn/TiXtzbYjt4F8AbZQOmNeHOBON/nBVM2ovQ7rxJZQ
r2i4h/YlwT4B4A4/uvrqmCLSK/ALwNier6nZP6VQPmx6JUaGtoOkwqL8g2YsG6/372V9Xoh4RTX+
e356gO8KdlmGIG3KnzxC8Py5rtwx2mAdYFswhq2+rzLM5oURDs4+lGymgzXSwfGdCZoJZlufpn7s
jW011SKWpeqT/Kmqh7TU4/yAReJ/dOwlHHDyLKfs4TCPsQH7q1/Euz+1l720vj9l4yPHILuvZcde
vlr4Op3DesaOZbhw/92C6KZLmVBCJso6VYjKQx0d+uSj0qs1Qk65BUs8Yxr08WvEsuS/1gV88reS
1OUMveB79YVRZgakZ1+2LQTCgSrehjZwJLMJulazkSwPTnpGADf9hQhOAe2uNE5Lgg1R555wkOB6
MLdAFLwFcjvnDy5vAmhAtZfvnTwwtyp9cAyedvpvQyuZeeUIH+/759OWxHdMxQEuMgN+iiztECE6
8mJttMkNR8G88pFcTz9DUFpVo5N/C/h8kX2d7RwTODUhcYQgjdeyi0bn0xvxDwD5f6UtAAnWptb/
GVV45sHE9DYz/A0KhfMshh25cw2gLr8ImDVLtEUYvNXa1eooCypyMh2v5pqJDFWGiwkZ2vvxeinH
zOzboVAkkcNd/jmRe3dB5KoTC9EaSi22AUCKgGhEFZs2/78o/NsJqfm5263JvWfUFO4N2BlQJw9z
ut9EAKL5/zdDOVtQ+wvTwPn9sckX0XOeW+LYMAtlEiXyfU9BfW5b7f5B1bSvHQeaNwb5Hy11BStW
YkkzIhdCwOxSq0s8gTSd85Kx1ixTzjsohiJR5dgTLWSvuk5AY5/HmryDw/ajtyLPPa2npXA/bzoP
yFnJH+oGaNJY1+vI3lpZ4CXwjrbKP5E7YEHg2HK5B0qLE9s4PvkfQrk828jNb9wPvG3fhG7JLU2e
uEfLAlX8XGaICt2H49fJeN+QcNIKQB/pr2wMqWwvqLmgqNhVZ6i4bBb0fKtQWOS/QyGYZN88gOBt
1Hq3K7mS4GNtVS9r+DK2ZsUQA2XmT8Vt34rUeVbi3dqClUPiATdAHT7wtnSGJCtGrGnxK4KoUj5x
/JeaGSDuDjzcUf/bvjG2lZuFoZGqeFrJ64E7FPBBmuc8INKjzGF3JkvffY9mEaaofGfQZKq1xI8g
Mi7VtoblhgMPOsMvslmVOBe091srpjOliVmP+jOqYPq+HiJoxTUCz9Rz4q7I4gQ9p26p8oNCzgYP
wAHPDPgvZZV5E4QRWtPbeok1av+iWeT8lpCsDYTJcIiLWzjfsg4SNvQ4aM6dkZYCH/zcxxqDIGAW
eUC7Jkq/wqE8uWtY4kFrZIcmmxwUYe/aTo8HurcOzskEliwjoV//wVEOzTBCuZakL8HU+sPdhKyU
5lvGbbTlS6baaFWB8Q0OHEQi2XrT5UdeV8LWTc0BFkfq0w/Vzl0V6DkHuj7SOsShnmuqAX+p3XRS
aEF31RdV/ZqoP9qYzw5yAH4UkCMAqLdPWKPfJ888r4GkNDxJj04tMCbajeIVVD61IDTMDzC7qfSL
KJotIj470eWTTDYdBNd8EiDvTfd/+mLjglgoCPF91YdCftj2YV3faqh8tLHczkoIkh9w/9mfB0Xd
cREnIFNoNYNGHpImtwda/X8+lo58a/Re+Hl1bsCry5/treZid4DspXEGF37DEpFwrpbY12TF/y8H
NHgg00k3/aTXA4kt5fnILZqGZ0QLuQzDMnFuxBhqRMIsBTKV0DNiUfTqh5PCBNfcy9xx45V4odEE
7mfPXiAKkah4Nnv5WW1XA71uVhhpDc8/zjQ8kDwnMqQYxPuVQ8CH47EhZgJWYuTi8TihmZJgd0Ga
V45p4z+zNUdqXFhkVjGYX0NPghAjQ9eFHGD/Q6cuwIyR0fiSSBPDslIVekeAh30jAFfXrXQFhDCP
TbPa80pimnjjIHDrtg52FxvBid07fAyzHYAbhGJFdAOPg/63uZtP0QINaBDOf8wlwubbAmT+fm3l
x3K8WCOe1ioYI4pvguJUwYXmcBsS6q9SD/zyX5gEFBza+3TToFIP2uR4czT/ZXJRl1DIEIOw1IWt
6Wc2mRdSCniTzPUzSz5i6BXtHdqodWgthYyYqV/578KIxM5+zpHaEv/2elTEmv5EbJ+1oPbJzmL0
cO+B6gHLFVQI0XrtGkiNDl1ZMLu0bbuvBduiX9THbySu6XT1sDcmR/TMqEVyQ6oHXg/L2Az0FQnX
JNk7PF9Ma6MWQXMPi2+M0I12/uHUOFX/kujikiC8M3pi62Xs8I4ksjNcQPohdTe/jfOIM8x1f8fB
M7Stl8WqCd/vxIkIOdiNqoSWQ5t4paQlgCyenwyK9ugtbO7d6Ex+B3dN5bu6AS2cqpypIKoDlBl+
U/GrStB2hPwXa00OD0jeEdkgcXnQFLlr1VgB+lZlkMygoolrZ7vRQNUlEyPYtY3V2GHqCpHYOg/q
5e2phYxDjQLrktm83V5aJKmBDn3uiv437oiWFH4m7Vj8OTAlEb9t1ALGw3cbTY1YSzCuFyJa+9+e
L99B8M1uHPfO+cfDK+7nRZC4xx9n5aIOoAuqgBdGAW/s73s8QLoW9wvQmvWh7LnDmRtYkANn/p0/
EAsqG399fJ+sat32IdmlPrqGW2QmejJHWqonA0biMMixXVJaX1Rr4UarI1oWnU5nHgVS7l7Ivqxp
55PVlkQb0r3wgFbGixT3gScYR3dSlqfNt2MEdVSILF7Z2/K3ji03sj44qLleb5QiUI02NKzN9Tv/
gaAyc7eCH7BHULiHUw0nHH8Kq8VGJwOy1CJukHnm7uvV6I5I1WZLGlWuMtk0wgWukWZYSHY/GkXr
+9fGDygC29vjEn1TOTWGuBO7NvZvGxgnz7ApOMTd9gG6WgGrbbtfz5Y1SxeDkH/Hn2X4JkuXzTvh
l1N90wR04O0y3JXv2OPy4MkMmzOI9E++GzUI0d58ZmyQJpQKtIL+oEQusTx2DNG2srUNfMW5k8Lm
29N1fxYQaoOEKD2jPYVZrSApUINNlcJ1cnm2uXLnE51FCffF8f8pt0FD+/GvqDt5m6Ikmkc0g6kQ
mjYUs3rn1zy+DYToxjfUYLV37T0vFrHVPNNZhypvVATKDJ+HwpyEhjd5JuMDa+S9+aJhdGvvuYfk
BcNxtjP9HkLGwwbVolNKdn5VlSVK5A6aFG5sJRm9+U/uMRshwIlrkcti8dDw1NTlR8UuIH31t8/G
z5NXssgMNW0ODVcUnPR24xr9pZQvhfehI1UoD88naFcDvO+bZeYxqU0V016wjeRWyxkgu0ePamTq
BeRUY6PSG/8dSwMIhM8dWkesy7pqo6Aup8mctyCdD86YteuCsuX98gRNsoq86XmjxdgteGjrJE2U
XNQ4S0h3SzJVNcSRHMQkzrS9CJ999xPsb6YISUK8Yg2hSRxojSGWZGnnunjEmyDOSDkzcufzSqE3
5H+eP0l3dwVgnjiDKmw5vRmh/Rjdx/dQ5URXPCRiUrnFFFYB0sY3EZ5muujCdPTylaJ8g2LbBLsL
ZSshqcaTOYhICL1/YEQpiN0IZlfSXRxYbx4LR+I9HIwf7o3eeq9XH06NEc/JkzdAz/jHXQ9ruJJa
YoNLKuezaWFkW6lQ7AnIlSAntshbkyWPMipkOdJI/OMFlSh5+Jj8qPkUHllBbMQ3xrJmkgM4qc/J
TUKVFvJfa3KZ9SHNzSe4FZr8onddP/S/JufGOfo87gi/NKqL9giBYUPiCBSGCCpMGA71ur0oRdxX
CBfn56NITeXuzalj1QULa3f7x+VTkNaiBdPagfNZVl3pwwur5mdlWgNZP3Ci34x1A5r9uBCKzs5C
yaXxJRCcMryDJa65BnXfAt6N9A1wfOOPeM7FKGZdbhuiJQdjt7/moBtsx+rmIeN8f+5tdDe6nnME
hs/CDRntg3CCiMqtQboh4EGL8g2nUoxxTlK/DSQnHodOG04rtpz7RvvM8JKpdrzkEtuW2G5cjBuQ
0QbssDKslkTHrhnZ0eRTboJmEEJpgcjoAfvA3snCdf3YERZ1Njg3t6CTcA18LQSIqPsLIIp5rU6W
nM7NAUAvf8dw3Q6hjLdRD/jo6evlYJPKBimMSsykbtLQq5W0eAjAIzn8LaMal2UH8dyhOwwea7g0
rP0HwyXcxwiSAWx8KiQbUgINRcXSsYYdxrWtQ2HvjeHzUbyX/8aEJQNbpwJUE/6i3vUapgkS6PLx
JJFhzoC855oXMJ4J4rSVGpVhgxAs5802ntYbRc1Ud/CWK1keZGYy8BxEzFmhwoujWiNdBm7tSOid
i0MCkwXhflfqLgOAZprizED94ckUDaPt12cwn3Vr38YrWZ9sSe4zsuz/JVsWOI3rD+EfC38BzHsU
FrPByl08kVFKbRm0+kT9lNBWaqGFegN/5mYjrNZTLFI3rC/l+20V+M0s2dyxfpx1Js5rLX0U/14j
eVonbfeKSwU1dOkjDIIA/JCe3s8DQVfpguKTMZHDpgS4Do0/QRJM5X08MW4w8RVIPpik2lFRD9lt
lXGT5j1jHW6NAYcTSG0tuPVai+VsK6phxfu6S0EBzT8d+lugAx5N6GYluSmc1/ZXF8qjFjvLG1fX
cZdVFTSMEmEArV3VcG2R7M9Ox4ObwZ527LenA+lecwF3UuCcSRdYEIAYJp2CYWjoQcEg7pwXiKVG
drFTtxN1ls1tOGU3IBXZ9NyF6e7hY+I+kMf1Myby7g4Kbd1BTlWI5perLJHG5VlwKyjP5/ZMgDDS
JpyOBIycqQoMcfV2BpcZu5F2tTra+ZnvIG2w9f3iJYZ3djNVrvfyAfMYF9oX40qyqrRil1mPOzuI
UJZzR3qlcPbDPp5QpT5JH+7qUy84fT7GB2gHYKuek/XwWabyKip7UQEOM/oaOGKtMHK5wuhf6Lx/
mdDzxxCZL5/4c78GET5Pw6JixgUGuNVdZUG1wDRGCX91EfRniQHHTB5DEQZ1Hsq4piaHcyk/RGEs
ROLSsRyIf7dJUiObbWqhTql2g0i5b2NR2DliI+oAu51BuMb6kr3jtDKuu9lcA/gmf6wQc3Q8RPCh
4oPEh1gJvnFYG28Tcu0mlabDjWn5EDBzV64eXPBD/DZgrM+qbr4xOBIIRRPSKHfiiDrngEBADWx9
/z4dctWXPk16EFOHnb+1BKxvCdJZcEKq3/UrgUM9oNaYPpGn6JZI46cEkwkKl858Qj3c8/0sJS1j
elW/kxhStHIfiEelFla8q2xfAbv1NuVrX5wfuQASPTyRhIr24gbnhShsEJnnFx2Zlp4C6vRcUa4W
nr5fEVbdXphA3bn37+EvdqC2xZmWR05B7h5kxlilS4sSPL7HOo55NpSrpUCjwuSyfvbELEZU4ZHB
xjpG9adgBqh0N07M6NaeyFsNloZYE8+21cojT0bRpKy3Km53ujw73LtePbqUh6jOmA0OuKBG+GtN
mohfSIqoZ3zmNU+kLN7nls5w2RW0fUYc2j22oFL5REvIfOBGyCkBqxRvE7hWYx1DYMc272VstDpg
rXlxWmANRHLz+du6IlyDadzHTMe42tPksNfR+xsKSr03dU05YeHO4iNPCPDGv04rPJdZfWNpLyKV
/EPJZiJwDyhqkkWWOq6leCwZKPGk37AyAyy72XjVrmllQhlU6RK193Z3ISk7uK+zTfbKigHI9s0N
oeKp/ltFRpFdRiKVC4oGmuDVQtZDziAajWXOzM6H+CA240hd1eIGUu5W99ul8+rruUtPW8tuD9AZ
ASXHastGrEXX6ri9GqLYNjVO5Yk9pSDcGjF9L2sERZaoUfD7YM3NsNxFH/GZW+SXMP2A6wGkjwss
qEEUAOr5u9F2ZP9aLrYxM4dn/Of6jkPwKmpAu0A0aVU+FQC8RmsHLcGkVUJ2bm2vhw50DPyZUokW
Qny0hPXkL9S1TZlBSPHrx7T5ojiJNWOsqHgHjHSU9auGloNBCPG8gBEe6eUMPUSAI4HAK/WN8dRA
H+RxVtOnrnT8fXdG/XlCVBwAzdNjievEx7IxaE7h5St4Pv0QBLaycNClns89zrbtbWRKqbwFRRcZ
BUaryAmP0Kb/T3dRZBeSJgVX3npzVZRZESoV72S5/BVtriOJJ/yN/s8ZYBGnHSe3JtRvsj3pE+if
dCSeQgLv2wrXoY2oepA78T1VXBp6dT/PEpL9zU6WEUNJxG6HCOqT7Tci4Zmo2si+89ZlpgLMK136
qew/gl5KSh8s5Dw/fWz/7qQlc+nV2d6QoSF7i8PSs/KC13YYhB2SlC5SOGvFJEMljsVS+QBhHBwN
fZ8kTK60hdhmdw3if64walaz09kFrqpSv2Mdl3D1lvSdbhZyebIdsyPjSYyM/TpJsn8YF/Yg9J05
Rm20eogoxCLP/uoIAULHKFVnLzax8qPsaWcU8qz7/qeUm+F2LKMyVVFzXJwhJ/XXuy3HkxDJ2ULM
jVTzLXQogWeSUVGFmCLoStYPjwPn2QdyEYnFRk6PfXTSVCehtjdsAw/Jdp585XjwimQm15SJafXn
Vxztixkup4nP/+60q7F9i9rmPZCEFdEG6EzQgRPTq5lnpsW5bKgu/9XNdxA8tamGvoly1Mct5sj3
UM9LPhrXUsLlT9sM7cvoWPmVRurb+DYJNxoN/vlSo5Eiv9cRRz96X8RpuMWA+OlTg/f74092WI8C
Vq+fxV/63HrR/rOazM3/VACFDDs8JELQriQn4rEBZEmADU3PseRyrGLVXqEykTFkUuemxbsWVyb/
oiFljC5YnDrB575YudiPmtFZqaIqZItti86TGE4XYWxunFC5PpGe7UPnaawJgVn7TJ4p4STkoTeA
VZ9TGAyaFgorTCKsIqJ/w9eJ02nZgjcwy31gkZIYj5d2jL1BFbi2IleZ/Y+wMlPy9l8MrRoFPWUZ
MljwF4Xs80I5DTIEOoM2TVAK/NZb0o3bULXVW+/Kb41bUajm5Xh58ensssG1Xf29Ras6XUEa+nO0
dJySOTXyYdTVd/HbtcrLlsjXVj5lVodGluG75ffaXYZSRBWJw0U3X8E1U8EF/59SPbKXu0pPxAfv
E9DXelBVwib0prLvcXycZwrVj+gyGUfbisq52wNyxopbAI6XuC4aMQv4ZMaGCf1EjFu46CM1uGSc
lrwpxmoMLPUIF4B8btP0BfBwuYx25hUEEB1b9GYiwIw6B+2rBtaA7tzdDYFXVifdKjb2IZ2Y7YTu
lKS79lp0EWq6f/3g9or3AeUKgMWrFoFRj2E/HsrQRTJBS3Ir+2m7pWQozo/dQzY+F/Yzs+ImBJ4h
eMg4kUKYAyPrLQj7WhUiEn8eRE7sTdB58IdyQfuIL292qN1o6Qwr+ZAz+IeNKS6Hxt1NHSuaoq81
+bHH3LG/IkanxCR6zD4fh5ozNGBvp6q1XHDTbd4OJyYfEEvqRL7fg5Luii7gJidEQaodjONLCape
KN8fqe8luy4BbKfRbbU6DbtwT+p6J2pjazUfRSfxYCDOoXMaWHkrn79/RR2AQhjzjvOX60XXfXKN
4I0TTIiFmhSBlNc46hCGwVV/RLBcHzulOzSKXl0woQdlOTT3qIYFYdYVKM+hjugg6sTcgLbIjdXK
hyHfDYJt5yYbzKnqwPTSSBFpa6dprPEVj5XYqxfpya37nQFm08ZYAYcw9oPITQdBz/tuUgJHMrjN
+oao01zbr6nvY4Mfqg+7kq2BO7UjG8/7IDQhp2bn+gBgjKSpkZBZPRN5hDl5KnKnrDck5kb2Rl3u
P1WlpTlUAFgUugkwhXKc3Ib2DUeXJPY3rxQgnU0XwDRCpgCAuRqGA0q8SHWxwTH70VXisJkcuOFO
qkvQgWCVkknqCMdJQxuMB2fhSap4JG9zimY1i4iUmzl/FPeN0Gg0x7bcefTBr32uqcejIxdTmxB6
8ZK5tHq0a+dT8O3A+jSHBUwspf4vt6jbF+j9YSxYzh4g8DSp038ObjilWI05+QG9KxqFA0ERU3Lx
kDFgCHX3JGKftFwRS/DZAwJpCskFFZZYuwt+hU8U0M+isTPpnVSp4QRMLwXOxuwY3wYT5JmalMcB
My7tL7dLPkbgbNcOyUbBO180CUTXCJRhPpHKFGDTaQfXsu/10EHclXYKeFEvRozenUAdsD0KY047
LNlEBR+tDSIkQFqjGDFlDcvb7hou/5p9xXzx2eWHQthcb0D1ysIgTbjgI63rntThRoWwm4BO0ln3
Pxh2RB1a9asjpeaw/buUHrVhKIygXyoJXHKYcW6doiaVpCpcz/dEIzSSW2S5NFrYXujDqBoURlgG
/0ZOGl7b/ugI1BGpTi84LNsSswD8vX+GitCAxOGkUzqenJvBESwjvrphdwfveoYkr+Mg/+FoBv+L
hpDSUZVwPNBnPcU2l9AU8fZ3uYXhL+5SM9vqvuLtd3bbJDXUGwzGtWvvKhXC/YT/MERUIxyToXip
EWuvlVP/zbztQxqNDxn/EPiHNx2bQKtjtAwuNKAQR0JDxeO8Ola3CGzA1+CT/rO8zza4uXnBdo95
XS1Gb+8Bg0OCYI08H8GwF44z5lJW00HntAtSa2x2u7XlEmRjW1fP6wcZYcF9erNOY5paCBzmsLUF
GfFNF5una7Bwq/3N+UVH10HMA2yCndE++QJRVNQC2+8wpDuf5r9pfPmaZ9YgKIhQL5cLiAj16KvB
uPZJq9sNWRmzCR3eIx5mYWJr8dFT0cU6YKKIlCHMiMWP7ZMvc68zcG587hx2NvMLV0nzv03gf0tK
5UTRp5RueVuJ+cZ4op3i3YMf6qaRjZAxMzS9FWt3XAZ+9q0mGeyC44N4GTtPn6ymO0c2hobSvVP5
15nzBq/HdlKAUKAE4XUj/L6RAKkL7sdmkGAqEVojzD4qBN8SfC85jsWmuP0D2sM09a+CF/eAV4Hr
5xeIO2szM4DeHtb2FhgSPRc9pHg68PN3V57xsDeZZHVywvyX6Ph14PTvd+2zDOeZNxjdJEzkReE8
tUbsPcRWsifxWONpwu5YFHuKH1Ag9tecvJ+H4B0wVPbxuvGzhitcKRD/ZWXqnDZaF7anS7j049QN
P4VGFTj5LFVeaFafjwct9rYlgtU6b4AZaAG3lBOMG6dcC6RWXMwZ4c8h/xgYvWGU98lMuDJNWmig
ToQ7HKIwITnp0wmUIczPDmkxRoVb3iBUqE8EkLFFiOxEl6p7fciT7W3k8avLg1svBwLv00Bn4rBZ
BUPffVJkp+OgL4eccC07wgnnFnP2MF3Ra9vxR9dSxKtSwIosi+N9+UD/r2iMRuNto+Yvs9+a/gle
vA7leaZQM2kIFQzJe9IlQVHBQinKoLC/J42Oee3eafffBoa6CSWhpSP4uXXMOKLaLZttZrA6vCrX
MHqSNxNbTUwFrmFuDlawQJkg0d6IKiC0K/oKg0GWKgGWanTlPBCouhlQoibN478mlrvMi9fAt1Wn
qKquWHNm5aSY9qJBTo1mUBqUUYenVAEdupfsoqFTPl+lCLLJQDQkFFjyW997eM+KZkVY38qPpPnJ
UnE6Wj7lW3LZojbcjExjQOA22QXa+Nv4iayNW7BLJwnaQwYyuep7JCdUvy9Cg9nub5yhKGkst2qm
Aj3t6ZHNbRzJpmkM27QRzR/GOYsEzlWWN67MuGtT/CDeL9ISFaBGzI3q7+tY5BRIUYOT+zYuMTqy
oD1gTkv6qZbeTiYPKqlGM5UatjnIeDy5zgN5rNuPoWkRKbNjybRqGFVMosLNjvEoQqqKLjkiO8Cx
UehKn7YkaOCjh9SSzGYshacvHM/8pBrrMD5n7mx4ZcmbqRoQG5mN0fgWGgohE2QFX8JBfa0X0L3z
ff5UDDx8fs8NLNe7FeT8RlgZlOQDBvff0ZYOE5+AmnOyqpBodhF9n8QdJXS23WetKvhHOiGlMTu2
gcgglbOCiG3ObyjsbryckDFsFpf+e63r+/6seLamosY3ucwX00vPTJtsrLinOI3xHQ1UH8FB8lbl
frirRSnoAVcP59Pawuuymp7DIOT8wEkIL84/fPJ35b/EEPySoN0jXJ8Zmp3STfwSD4JWgS72dwFx
bDANAgXTOWsDVZ5tgdUlel7BZNLZ6Gf8AW10SoQy0+6bEUTSYBR7vDr376klzo+KBh2YztgRZbWl
326nEcrGFzTPR+q0IwASFstYehvnuwXYnFwA393FbH9eIUZaEOuO1OEZSw5Q8kCeEZtNbSdhh8Hr
yk9T24yEc08tWlCpS+825G/oOhCJPGo1EA8n3rSSnV3CyP01RtuTIhLTobiGg194aPery1gyog5f
438jkkTe30sza/WFGbGT/q4Se9+mUC6oB7IekR0kqXjk6qGNUQjttAzH5Fdy4eM2KEMEKtRaJc1j
rMNMbx0MK9RUgbwyuy9ie3LHGX0dAMiR2KLFd32mSTVgPuNNqg5pqTbV6ykPy8oIxhL4aJcjlOaz
DsBuQxr/hthyZhWeMoX0CzbL8mnKbW48G9ZuFxku+gT4k2GjPHPzxRDXUFtU3DmQbLEttDRseTKj
PhhLGNCSU5wPL5iYmjdNyfrb1eBiFWXLK6I1iXjsgXK75qcmmBcYjzv/132aLBELZgRyva89YHJF
Q4bLTB36InLZ3yMPuDKX0CWWXafzIJhFgWbGViE9nAwfshYHLDordKNH38Na+Fb+NRwquD4MGYHb
ktc65TpsDj0MTcuWc5dbVMWwPOf2VuXnCtpxnT/CZOiXmJuYA2lT/Hx5LGam4cTwwL1Yz4hr3aOn
6fsL1psKN0wbzjV6TQur12DJczD9MsukoTIbkUYVkMwqPQ9IBPJM/j/C/U9F90YN3RhjdwDKeo+G
mt0sCDAg5yB20Fy9FOBnhsJUHt0JYW8qEIQlVjPKs/TaP9KztMtZ3twtRxlqTRYOMO/qugGSzzHk
fQEqTIHmdmKyrZ0f3r+v0eU4sjE53IMGQZlXCqr/zujw+bBnkQ7WyPx4ef19YCXxD678c/tvk5Qd
PHMRsCiGwCOh1jByIRrn7ddeM8FUWiNiJbGY/yDXwttix1Zzu3R/pOydIURnueh114GzW3EweboA
RGSKiy4sREdysHo5TN4+EqS5KBU78aEyebmXrln5tXho3PWARHpwEzklsLW3yBiFEgxPxjEyGwvu
/kKlDRYnMsymqY2HyZqMBOpnakIj41IDdL/DLGwo7NgyRBMFl4s2yuR07/GGyWrAdRP2W8toSQKt
PjseMIOBcZQHFsgj/WmuEpwgmqUftUiOsMDBQ3J9WfnGEhk36trAVoOtK8oPYhB7Tf9dzKYZRNhA
w33dsBfJCviW5M3WaZZB3zRsSFmhAmThqIhSUNvJj0S8elNSawS/kD1XO17fv6WTajkVN0vtSl8f
/gG+Gb4The36ek24kV7CPr+Mt1pEvD6JLnBQIP5F04TLDFzz4l6JGYH1gpzkBcCz23Izx1zfL+qs
C7FlfoMd04w1C2yPhjMqduPUHtrHUCZZxaUyU6n23vWTMJZWFhXuWvTuKebCoDWU9E94QJwaRIpg
8iKoRBuhSgAc3yJYXy/W6mHhkpRNu8gX+TYBFca7OkANDEgkN6kVl1VxMsRJBj0UOSA6QX+S2c38
ww/ECRvq3nLf7yX+WJuuhcACb/4+zuZTGQq2F3/LIKup9wYyzNxl8gctqiak1omZyOJimbkqYTmK
pbJ2g9rsH9qP8cJirn9YiDrBY65JP1W0Bo/iQeQszq2xWS8PruvVy8/48z80ZCV1oDJzaM4eZ0CN
vgXC8u0J2NeC5d1Dcdeq9G6TNuirUIpL7Fh3gvyq2MDtmettNAp6e1KeXJ9uZPkbsNbxQUque+k3
jk4VB14DJc5YF9etbm71Ni1smNREPuZ/kJoddGXLNIXpyHwlfjTnN49uDeKQmQk/vCOjliVKG8q5
9Jg5L1uE2sfq6og1qIBkg4l2CT9Hq3dYRvcpWpQTb2gCaRyz4tdmClMun073X6PN86XysxqaRxO5
LapEj7WXzcR5DTAPUx9JzY3uAk4Ag9lk0sJjRvkPozg3p4PeCVVWYf+vQXIf0I0RjuFfo96hm4Cu
4BBSkD/BZmqDYm71qoFDMizTths1o5fxwuXXrUZUUzlRCELypay+lgxshoWWAGVTjIi6ocEDNzfY
1sY5Sf9ZkEwXrVPnyZeEN3WzuCRHqHFfG9CQ81BMpYYl8PcdMgblayV7TTECjTUJy7k/UqgSWoR8
J/6aOPaAMIGAGjN/vYxtctGEjTKpleqE4IsZXPA7L/ue0jcCP5axomzOBiDqrQOWR4aHiVaE1apx
KpOjuqEWX0fKWfARXMcydQPCNHHu1bYViZet4bdY7lXwL4phRE9C5lznDRgRY5a1tAQd1uubwMYt
mOZc6wSbeRgC03Drnsph2RKGFYSNHT+QXggqVB9xMXKtEBvV3o/V2v90ekq7mjWOLMmpHVe333oH
xz+B3+AXGgRE5KJVjvNKc/97/YypffMeYHjMDn9NMZaaz+7fhg65lOWrOrXmiTjCOo32436dFQaE
yZqWaIKu6tBiILo01RnnPvGltaOmKWlyPuSnqjr3mtvq4sUtl990iBHmle3evgfsQ3GGi1TK3YR3
stAetF3v6rS3/yRUkgljzWnCyglPi8L/9uRe42Seu6QbaQewrfEESeZmAGaUnIzPap1c56dLjlyw
XE9qBAUggiwdsnOJAMQl9O07V6JHMmjCY4YMxG5UkTOBc6GHvalta/LES1/AE4quj75hdZ3Wq4jR
nPHpzoo3kJZQOFc0KNiA/3Rk4Q35QPWdtmcvDiOAs2y5ehmbl8VpxalZO01UkLsB2qmpQ4KslMBh
IRpb/ItN5DyGFsAG+c/fX/to0kgHtO2aeB6HaIKbn+OXXq52PDnIJR6hw0c2WJwk4zmoK5V4qEK6
gW61aj1HhE06aLzK4rK0Qgd/INZ4V/rw0RiFClhE2qzUplKb3xAaioVlAvpc+chzWzNloyarqDah
opmS6UxPNyrtR0Ce01+LNqa+5uSwEq3/CsLlOpq0yGZ4LVKwuUmFeq6hsnMQCunhR/zdzxzxLW3Y
Hi+2wG7hORaR0qNsEXaoWLScNRYTxK+8UOK38OaFuDF2mg3QbY8eGP4q09+m9PvRe85UxxvBFUhU
X5wRVH0TX26jVAD7HfMr/yekqU4f8kCcK4grvVAHgP89LiBtzRkKFTqSmSXq1gZ0Zq4wUs29y14c
iezGXwwzFZLGOhchA8LBtk+OhAiIZGUQxktQKG/maqAAnv9TW4+BTBgOlk4t3JpWU3noXrGj86Ot
eVXMH5WR4FL4SrR5p5GrYyc3ZtPPfs3KJvSh7NQ0hk+5IZR+ROqE/M9tLCrtW07GdRcOaQhtd2mU
5zQyQNOo5WuY2t2Q8aNIcR0+oed/+HgdYooqduHKsRSGC/Jhc0G+4ovSWRpGPXE6VGnOGBSsMWMQ
cvw5UJxSdiF/i7NAbBmRIcwKlxyEAYsoDEml66W0XjxvCRSMTNGHT4+xYBtm4jMtQQPpoPFVLRgH
i1x3JQdYp4dGbQmAKlmsswL6Ed82ijRHHp2zsclk1oie+LQULLUn2caff84LyKBdAOXtf9Ky6qvF
Of+QjNSj33/ylKwTJIE1DdkV0OhgPxagz/ggUo2XUtIn1Zj4YJVPLe7LOl6OZhHYrOhBAStMC3La
uClcKnGGwjiwNDczEHvN3nuZdj6SWF4cRZ33tQTgmWSim+Vjho8coKrd/x7kofviqCAJzZC+eT0A
ouqscf/L+UQMfIS6I1IOHl+uqwF7MLvqPkLieZ3unTSaBkOgqlQvHoK+ib2YCKUFHz1IzESxtrxD
l+zx6fG5g/rwZCqrpMwsCKHA5omiVpP566evpNpHndTyfzJAO1tYDkxwXyYWJYCQ9Gc9nVycrGO3
Rj598xGN5lDNRdie4LTtMVJLbL2lNKtSTAn4TSVlqVWr/24puhmdoaR2iBlRTPYop3H+aeZ4bDxU
HuqiZ+JBRyAgiZIX2TB+DG59+71i1wk9oBtQ9ltkzoTrz4VdxZVOD1Qe+WyTiNQjF2DXdYzJK5/N
89GmxgnC8gnwqTOZjtoCelN5O4Iss+3bztwKjs/kKQgY+pqEj49esauc30xdkDsAPOIPZ5UD9vNa
jeioArpD8Nt8Y0GspyNAJa8rOnhw6cP/G8ToFpvegvVol7g/0dfIMc3RolTlRo7jlhANEL++eTr9
7VWqG/DriIQAIZEk/4tdRAoU4LNVMJsdsRG3oZLjqr2sdDO82qwqj/Ri65JEvw4L0vYnppLlH571
4xil2ENkaeHF3lVXdL0DoUxDnfC+co7m4IC36kyGEpJ9xs6gx5rBiqy8iRd9zdw8o61cpQwIzNKg
kRIMOAm1BcJ01LWQWAyd8KNarspML+IGhvGBkwqkDdoX2HE4Cw2un09CNFcslu032dE+vxGeIbkV
h++79yMAdlC7EqFdtZhdj6Pg8REh4N4EjRZMwPPWVcLvrflC+2vsXKfqt3pK0PIUDnbP4D1Dq4q0
n/PWMzJWlcCbsOgy9lqR45u7ZPKDzbGGXM1fDl1tW1jh9d/FTS4hknr+ThJ8ubRjEidCGDVBHpPw
UFtDbG6ULBwf0bj2z8QSieMj+gyx/lsT+cpTmxOrTOmDe3ImmF9GmsySaYtQaTqWoOfJt+Oo0v8S
l4IHAwQdk2vAPocxWJ9vKPfjKzJs2A146Bqy+2ZVQorunTo6yJzlisgKjvd7vrFLko0imDGlGaQb
grH+ORwhr60N0S4dkajJpn9sd7zYDK1fqgohMipyKrdbKX0V15BFpgAr579SsY6IyxjAhyEWtq3v
svO5RpfrEqsTjDwnJvvj7fbpdymU5WqUHQvJh+hjT03Pyrxat/KcTajx1AJLb76YGcQyeq2ZuAmt
NzHr0f0048F7TkxXKFNwKEfOUPlURi9wFitH1jrDLQcujVZAklyiBuqz1Zg2+Okxx4iifvdxKx3q
fhthcY6GfuuZcLTxR5Ze34l5K9q6ua111CNYy1FvGoS2rm1e+BCXbIXyiEmI/S1bFtLcSyBVQTF7
OGdB8/KKtd9EvxcrojQ1JkNOXCYkTCHHLtxYgEM+rTj7T12Ikp7aWIsazB7abH/XcHMdsTlB3rRV
P7YLtmSvc+OdfbSujfPcZf1Z2ZbGv0MXg0vqIWPuaMkf5ODDOqC3l2taYLeC3OqAhRFaLvkW1U8E
cqECrRy4/AlaCZ35rMPy30bc35KhdfKv1vNsstpm8RmVsnWNzPRNoN2CG7eK8m3JFt5kdD1TZLMd
tquFsmUb9qWFMlOGmLrhTWv0rCZpR/Nw5ho8XfB98NNlw9X1xgNLxAmCzzZpwNOEOIbBX6+AHgs2
xRXm8A2mUirOgDedSab7nNaAoXL42J/UXueb1ASym+zqmU1qsBkExm0MASvNqSQAy0JSOcOmV3NL
kNUJDN9WMh609F6UF7B2uyFP+lQf+xxZWj6R6fNu1/mmx1Z3ttCTwWUu6iwGazMHcGObApsezg+V
DRBlULDEkPjByjwnFX8UTcchg4OpaQLjjPaIXOZz5BtNUFPw/5ol1lrW+7hewaqGJ8q8KuGMrN8o
NJYOC7xsROqnqkCbsEJdANMi8LgjSersPhiFaa9C58h/vU5Fyk+QV5ogkpB1vbDEAk3Rhf6z74Ze
gHlcbjHLJ8Ed6O+O/xpHGFrHuHvwaSIbD6zoRbVBDFZR48lobyLLrtecqni3I0HNfufVp0R5O7IO
FByhtf9C0bJI76jRIWD0Hoamd6mqmc5Zd4LVByu822OF1/YfrldsjpAMhZpu6nPFhURSULcrQ78R
HgVBQr8fF9KyU5w5P69NsL/au33E/PCFxGhiKpZDl2O56UpRIiGFzQfwNAiuES0cQihJdOIqin/h
3Bp1xD6kIqIEBL0T5NfEIh5OGGM2y82aHMLTU7vH2NUDhv3aFy2j4Mk3GY3IZarhhTsRCfYzxEyD
oOZCGg2jkTNWitgdoJOSEn3aOuZJpCfx7IhIxHdLWSgnlNaja+HTbx9yn4Y1EM5u1Shi/vQ1+anV
lwwgCUkmHfW3aeJyaFVOUgYtiT/JTcjhUrKj+KcEZWtgOX7EW4Z3tWXDRZLaIfmOFgvTLfNz5wVT
jJHyyAgulg5raNnaQIuIF3PXoXonO2rn0FQrSCweFCjWta4JNKzcjWc3NcaiPhhypD9Vg1CyWmQA
2FX1l49o6nL5+BmfPuwVJjRu9vmZdgTzKrKZminSOs3CrHDe1zn8gQCpqlzK0QZRr74mdLIIPUrH
4n/LSz4grWs0D7fZTndo59aq7gCLIXmT0zq+I37miVxwa8h+j9vH9hH8ni0weTJGk/RcP3FBkyv9
4iMDma0BQKImtVf1XYSWldHrBqjxiatGHIEWz0gzJr9ZVhe6WKfb0BB84QSXv0qGUTXCpNiwztt6
+7M1ifAHZYP16hyfC30aPknxtHTgtUJ1lRVFiuArNqXysxj7HyFNvLDKwTVbO0yWbwZmOFZy/0wN
WnkD7r/OpVfMOWB7TTjp4amA5s+WvNM/sQL0zWAwNSGEW5oNOfIEDm5I2XJe5bj+On7jYkwHjfJi
mw/LsWeoHselXGKXpHkffujK78c9QSdA139/FOODvuHPF+w84q1Ru1SrUkUBkMgoS/RbxgxheVaU
FW2mAps8XwAsX+Sa7akMIejbMrhstBka/JlH2MiHXXpQEuh0/4nexlj0RJhb1NI8Yg5IE3FRvgjV
DYgynq+7bkAzM82cE1abjLpb7RUITA/3e6+X+pu2T0kiExnruHNqVVXgGB892ogiGEqeEFmZP/SP
8OF11bfY0xhtSRsIOtd3SxyM3CEntWSpoD1NsjQANio5b64k9WID3JVSsggBJ+O8KTQ6zuLLBBA4
qF61yC+NnO7nVhk/8bx9iNg9qROS5P0adLxkG4CU1wU/93N2esTClvrVelImZxvftf20pB1AD3w6
Hs6L969sCTaoYijE0KpsA2LgAo3QyF15TKKblOwxvi2jJvP+oJKxsR0K2GwNktALFcU2oS77lU0a
TEnby/e7tahPZ+qfHbJ6qYyIdxkFtGGGFLODGM5z+dEKd5HT7acYMA9q4tEzBlv4DPIZP7jHvDZ+
1ZhRYEbdTAcvdGYTLyZ+s/xrzblLvjmHNtG9gOXUTPVte42ZvMRrTaKu4tVX2xlIa14tkCmminU9
yVIKZ/ClzNjOA503izMeeT5LpVTkJ/RYKw6zSJX+1qL7YwOSILbY6dffbZK8Eg688f8mRSzhizYX
XXVLxKBDjEXzAN8hOPWaVVJV4z+jXzKzvSS2pctHUf7/t69hABRNbFD+tfqEcWdbSAP4bMYoR2rG
rYQ9qbvs/K46O98sl8DtQUgXHTqepls9URLAZoJUc9g2uEL1RYFRprBzx0MKxw4e9HxU+m8cUQht
tCRnoQar/+149jkTBBzVPivoFSCcbf1tweIhcFSohDqD1nCENcBFsS6vKp3TilUxvcreD0+TdR22
tfjiTauS9YaDmILLeQDL5gaBxw/jifivdQeKWtISYZhfxQN1YhSyPpfTA3gcN5Pd1YgaRzZ6a9pt
NBV0jp/PixH0y+f9pcP28V3hy0geBxtR2rm4bgn3jHKZuWHkSiVoLmlJrZvzyHHfbd7ohnFFGYdV
6T5e5FzHMAVMSppn9BJXKjApvSo660ZNtMr4uUbEkeIbVVP31X/G4kPzHvc9+831ctqtdzZzgxZv
ZDoxuyBJHR1Y7FwiuPFvEzA5lhIz/+p6ZCsJ60BcnbPky9s6vPhCF7DszFTOE8YAs89pkTSJntVQ
TV2qZP1zkyXuRsf5MATo8D+C1eUlOt3tItxtaOWWtEefEzj3eyWte8mjnNY6KEKRI+tTlOSubQcj
4843lpU5BSbcrI7XAFNlbgIZ60QomnA6jcwgABnE+KcdDlkXahLyk4o45LEAN3/zM5t/1TAca7zh
/UFUNtCr+0K5c6fn24AD9mEQ2jleiuA9fuL9xk6h4FAckVZ8njFer1U9b9O5RZ+K/kBQ0u80ftxB
EIWY9cDCdCQNHQg3L+d4vZ0Fa1LYE7wuMHisMlknkoxKTmasB7G7GtcjqauzvrLENY8HHpkTcn2s
CwtPeCsjcH9kBP5r7QDsvy5TABJZWQ5J9LXWxuRqE77ksju5shjjy7g9n62qVnmzAFxA3LRwvlpO
A52PmZojdDyK87QZq7GoHeLr40+ZkLm0Gre26POcJQrnJhQtfmf96h5LNTt/faCiEO3E8Stihm/p
AG2xFV9CIzEctmAl5pEmGUAmKFUrY+9zVm64hTg1u0pKFH+P3SKckqCYmZBqqmfr/G3UCxU4MQtJ
xjP7WUAImtxn7ZQ9VLM3RZsOZRapKSDvthvfEcfeCN1H918oEyLwB15LFZcu7VlZj9Z/rPH5Ihcw
0mUit8YQDNyVAEJc+5piL0zt+I5mAvbWK+maY6lKrmkuJsHHf27gl6/brwB0dql5OlqTwYCjmmRu
xRE9c60cFTLH0KCVXakJ3EPuswzLKQA5b500FpvvSsAO8gPaJ86zICe6HY4Zl2hpBxupfQUFJUuD
1bf+LLOWG1guDBIQJ98RTRekQPMx2k3jX8ZFP7IM2utGBSi/BRL3AetSGsKZEilUJTc9wckjIcNx
EUb9BUssalMmpLi0BEUAn4cVI/ak8ZfsrWO/VVOiVNArRoCG8/DBC+VeycOT8eqtprApzznHnmjk
gWQcOIepGuPCIG6g490p1IQhz75zx/lSFXHxHdnaA25GO1LCTLA/3rl9x7mf5uuBU1zhREftSvz9
PXwfQWRg2moDpnwREiUtiB0UK2q96r/pSBP/XEQRbYk1myDIVl1T7OnwJ2U3OZ8pMVZOohKpNpDe
ekcWP5Kq+6CrCB31d9GrvPOD3GaJ2BYMfjqNwVLUgrpme0IFU5DI7R72Trzcf/gunn3TKndVF7H2
prjNRmfp4uRyzxoJRxLH5ljUkbsRfqtiW8Q9C3Tve2U/08YIveQhql4Iz15ow7kwOLZ2ptCZ+C4A
Aq1vczY0qUlL6d0/HowvfUrMAlVzGHTz/FZWI645aGKYBYocpB/pFMajIZU7CXhJXN974el/R2GO
vxm3PN31Tgti1GCQGQFsszcRwmF6oKfB4SXxQq21CvKM/YR/B47evpenXgWpevLjtHvJ33ktQetM
Eh35SGYDvKYtuDCY5WZgnway9+FGX6DmYJVMx5qjbdcxqd9ASUEmGmLogEdYJpuu1Cqka2Yf6WkX
xyegDlti8oX2WnSFHzVW+zfdkm7XYx5N/QhiS6eHpGKLMe1x/y0V2H+WWOL3qJ0uMCWrvkSg+G04
US+EZKm5nKsvOYWuwrRMECHVJjjfzMi9k6vKlqVX/p3pHzSHckZ/C/5oR6c2ZT5xpolFIuzwDfQd
hXTepIySxOTwjrCyTys9pUlIyf2FssyuoUUYlCu1pB1F/9FDDytEd8QY72k91GWXU+t4gCjpTLKa
6aEkir+OWlH5Q7u0nF7MdsG+gA0QN75TD20rzXs4dIqNhxgoPqyFiqzi4CtpIKVGVuPHLRApuS5h
MYusmmFGY0h+LRiAdgIKZKCUCsXC7IxmaZEx7bWeqI87up5XvOkNNpuRnqI2/EIgQ5NKXcFRn75G
SVgtX65FGD0M6WLXGU4BtFE0xrbyS2vrniMxOncanp66HSU2OGx9nlXCmXhzSc4FOiD3r24qMh+i
kovqDi2STwmK4Q2cKWsKq/40Zf3a3GGswReJOmld8S9FEKzf7MxmXonk3y+fm13f1WQ2S+qBwifq
5n94Yf1OpS4hh4sTCPrZ7AF/2tlJ1wK+Gwl7xY1v+P8w1OmQ/XJV95SV79sy5eFWO++hiVhbCeiq
yGwmslDnRLCPTB82EA5CNeCDh5x+UX6nPhdtGT3uvWyWl/XnhYquw1G0Bsijl9ex2+9hN69oF5LX
m/S88QemclPa1ZDHT6jBVBY2naT4vBsuV8EmasZdQkXF05k66oDpQG8Awb4rx0enFjpw5PgbeUNy
3Q9hHmdaRy8XMGHxZUOMbA1KmjqgF4JheAgJwBfa7P2FrCKFnv6uYEbWcpgP20moil0UD1Y9ZdeO
JstwqTIVMFbg/9LpCferN/5lPV+vHszmDRueawc4PIRXlkh9k2pbMB7rpVvKNONOqvNjqcBmDHs/
KzkOwcHfrA9LkGNhfQ+18onItggu956lziHQv5BAeWiAVL3TptJTM2bXZISrwyHkxkV+lO3h++3w
oUNbfyMhgjNK1kliS8tFNEZtloqmm47jKs8mJ1BMYYI667Df99uA8Jap2+3wu0x9wWLC9Va/ibE5
nYLeA8dya0G8ypFb6JbjZmaBaMkrQ2qcvWTWBgfP9mgPXMTzEYdMOEIU1DGNCGmwQsg6TvBRc0aB
VZ2dPovsSERh4M3EjryjV9ACm7SI5kR5gsBGW0b6n9D3qUokS5QgXejXV/s7rk35/nX/VMTiKt0g
dNy9HmlrCxaOvXr7TrDc7S8pHc18bY38lC3zsT/TBHfOsExadsdhT+GInahbSEeOg8bHdxIO7bOk
Yegrp7U7zPxB5ZZLOUk0geAFNr9rvzKHLEQUM5b245YJ6quJ/wtSU+qQ1GS/B1oUDeW8gdjcFJ1x
cVLqDhqL/EF9S1RaN/tMzpckoDFOomb8d67ypmT4FsYLIYKRRmez4dhcmvE/kUD+PQa6iqBhtg4i
xNTl0OYQTaYDhfwj7a4GXekDjHbKHMPATUbHtwPX5sZjVE7sgfdFDu3FpjyGS2crPitX9kStByW1
PawLUy3a/4CjczZl2WhxMZ7HvQUmt5rd9wB2TZAT2D3IF26Wssq0KLyje3Nxmm+/PosPm6ODDaDR
yaeIP/3FXKK4iYu2zMU2OyS0QZa1I3+oIvfDLSUpUuJQZkyb8CxYdX6sn4V4m7CAAvIsR6vZR3Ig
aaSGYDYt5kz3FFuOAzOuR1o3ke8Vb+bQxFi9BxLdzv5aKY9nU+kT/aJq18zUKsph+mFnTFps5a3k
Cqx/hkQ3NH5wccWVYs90ZZQM8nLWzEUl5eKqcOGSHv/BAiO2PZxI/nhzsGFaftxse87S4EzXLxUW
X4YzNGVuzPCeFPZJmRYw2px6QbSPxvbyqal2B5q0ttaqbgTsI0vFxMjuhVOIeNW9qCPtJRf4cAH+
ekzTZ5ABPORU7PFuDq4NmXpVvtDw9XYOdWenOnB4ShSfgk1pTX/59mR71kFQDA29Zy1oxzFuEJ+6
JH6FhO4bqtySdSOeot6FOiaJUktIphidMxzIDH1kpqCtzhulNVn57MlmgHbUzt+NuOLPmF1r5T7+
PC/pp2UaFsyR5XkHHszu73nrrvdbo/Xa9BXEX+QoSQM4dpjfvmgNLXHZvcHeYl6rI48O4i0yUecK
fHm4zlI+ZZQ6/ahA4iq/uSPLPD4mKeNdCZP0TUM8E7v8nC9IZxcaC/L5DNlUfKGNsChrjgyZbcof
/rrIJVNUtwxkHLmcyuFQRw+mK9KuDjci1R6zohUhR+xfatl0c9AYjE2aMh/2p6nLLQnw8yL6A+za
Ui2DDcBAPyQyZ0Ikk0YHJzFFZA/GrHNxjnpS8hmdtUF8v8Qkfk7Ivy26Ml3ym1GXSabsNT6ax27G
quA0ImHx1FFN0X6aPsGbPhljx/nxG0j8QcRAbjl3ecl32Boxz28f4gVjiu7j8fgCtFhypSM4r2Y2
u7BOEFKfII1WQq4K1D3CcVP5Teo0CL9aQuZlhdOJ3nOE2Xq9rIJRoHlWmOY+8eY7VG2p2MqwT5LS
5BotpZb0sC1ZtYsUe1Qld1aJb2KWOzaRaR/meDpdjTSy6k+ssJkhlgVyEUJl2yZ56fMoRG7r4BvQ
+/gzuO/mf56QC/zIoUcmSAZUbBavr51jL9LnNvbukpkF91rDJmG77gsjKLiKiK0FGlCChzLmJcuB
eD5XERY21O64n+WH+rTCppCNp9rYNvaif5c1eIfRg3SGaTPzRFjhdvpRsq/HbGZeo7gc0In8IVsv
vaVMk5sipif2ixN10qUSZAIsGPAOCtLIxobEE3qnTdC8OpAJZl/8QcJs5WoxZ1PR3PdvJ76G3YuZ
FANHXrRegFjDrylX8GM1KiqAE3N8M6UaUB4SiyFyBZwRiUQZa8sVLD78kJVbR7FU/Bc1jQP9g/j8
7HN2DfOCueSOjmSGGkiVCeluefPwxRS6W5Yq4TRTNLxDdsKrRGuGSufaHYln9Dzqm0VK7H3ctNeG
jrArjMFAxyUyK/Qpm+LYBoYvEXAfxgXK5qclpwQgiKHadYFBAIUX7I2yTosYsQyfL2pH4k9L1g6f
1KtAEV/I/rU7qNZHGLo3PZdG4p9rGWC9o7fj1DjgBYIAgUHHCSDH87MjIw2BtXZfyFPVSIjbleLL
COU6j5WDyzZmZFuD0lK475uDDSJxEk16sA6CJHn8zWKhOAnE4xw3I9Ng4370xMnXShoLs/uw1Nz2
10ccmuoboykz1BvQAkpqz5yi+KFSS9b1t22QSuKPrhpYW/Ujgeu0vqYcBcF4fvx0D+0AYXBm+BTH
mDc13laIUQK1Aqaub9Kx+F9oM1LWgdwxQuwgMXqWF5mASMeZQXKHEdxqYhEgXpKcSYFmim3iQSW1
jsaPsYUG1gHgRp1ngwBGxvbCQNOGRc5uPnq2bbv5Md0HvfbMaF+SHfpiDh7BI53bqNk2i6eGFDgT
lT/RyxhVznSxst2rrtE7nSmpvCNaTPW9VQX+PQuU0jrfbAN/1YeXnJzvQeBpm1bGtrcyIZENenQc
dNeZ6tJWWwKARGCsWKg7prr+ad2Cznqadtw7e3e1qZYlbWWQmJCrYp6gy9sXlWcd+StEPQVK9+7m
hOl4DKQP1wVeKUX2rEeE7Y5MjYxPq23l7x6wIRw/O8LKtauAmj0UgC4dhdCYi2bvQqiTof75mmgM
fC3K6GZmmxMrR4kVukWB30ZUfXBiCzwKzXsm92PQh6S3FqWmaxKSAAxWsoOAj5K9fFijjIH5WSwz
iIkFc33iKC62uBWmHmIcletLdrJINaP/rIlmiLmicoq0Fgcsitpvv4G7f71YUT72jgapPEmGe6Py
rZ81iOVcqzllYJvhuUV4F0qxPd8F1ETwo4xduZoEHo0988AsTHQDGOO6P/fFjxxd/pHTw344U6xc
7p905it6QzE+iG4ExBQwwd6OCEsaFrk2RbCha3CVp61hpLLvFYmUmDo7K77isvIlX5KldgTL3TRg
FOPZObFsP//edhpCTUrb4yg88N7R1e0fgo6Gnx1GvRBopriSA8G1mQ8Gg8kFkefOGdw2juuqCIGt
6gA4JHeY6g8XhCG1VuURnbHGBbWpu5KbgZgHEdc/KN7m13vn97PPDMldhYxdTKiusooja6sc7DKz
WrqMM7lr542zOiFUjclkI7E0JTfh+Iw7aorB3Np6e4LwVTsncgZpHcvnUi19ABXBNslejx3FlvQe
4fCVCPCkbQJmWfQKXgC2+EwHURb5eXli4C0PlLRYzVzDoa2sFqdEg3erBJ4Hi3971NoR88MWgCAU
Lsfx6ilkZhT+6IYnYlnJvp+mRNQ3yjdEMkORc0O1Ng55LVa7faw2kdJFfdpd7WkPZaSxagF/6Du4
ipOK2FYIfjI7JD1cDM9ibgJbJEurCUUPTlqIKOBCLcU9CeEBqb7EF1V5OnCNLC+HbFHk51LEeU0/
h/gMcVDfJLLVim9P0u+kdHaJoqTzCKW351913i182lJfC6HdYlLD3Z/MhOK28vmWsUYocP1omRB6
pJiWpoGOfj1dYOxBVpw6pbHWdhZUp0ZlNRt3g08kC76v5lWFV0p9TsztBjVk0EauvTHmKagL2E4S
Hq8cQVGSwPWBEFQTubCn3pVT+sfx6D0Q14ykHOJ5zAKpbj3/hh2LqsDRVIgcLPHWGU8qGhUnGmYf
YbnwrY7yAkVIfu9Boa/HAHiMLNnJIgxMFjLbzmKyHrsQ4HQP8ux9GIz6Fl/77K1OZcIWBnFleA6x
mMHVN20e+t994VWdj6iss2otTzRYuzxdOPRFlls87LzpUE2R2KVZ8iFqciiADpnvezkVC4KH2Mv8
BKisoIvvhUWrGjd+T0LKklr9JrMzIkbRwIKtyJFqkEzvTNwkYLX3JqaM9qh9UbM6+DlbWNnQ7KDs
kJ7arBZnYK3pbFCBSsnBYrzIIKHi6w2BridyMyYxse/B2vQ/A03GtGft+4VNz1sBMdYw78g+aiMH
YeglUkq5tJqr1dky9DniQclJTfWLNNnHYhHPL4uSFlMQNL/uuoKNQwODxZgm9Tp4ybKWhklDKGJ3
slLsx9MbdoppkIuKhfPuSu91gfz2wAVR0/ecAp7pYGm3z+7XlTtv+U520XtIVsHzSRsBTRlumdod
VvModyoI6LPe6YevtfQtIEgNDWMG7sMJInx+6j5TyJsXTKe63EilNZoRIKCYXZS5MB7eVfE5E7pC
XNzs7+2QEkrljvKHOPPe0gWcuGDjAgYSKqIUqlnFQr/mCrhm4gxtyirHp23PP13NAmXg6EiLJmDe
wk9ymclGiMJj3JuD9AyRedHHuJtffIO1+wWdh6q8xUk+OFk/Kk7vc8hbQTLohMc7dDiNeQlwwvKm
28eLuvjdOG1xbC+veFn2TaE+x03HaDrvGRVLHDq8qN1MjAwUee5ydjev4WQnNNCFXAWlCwLrQDxx
+fA8dyi1SqtO7e/rX6lB2ADF9DiGVwaj2rpQ9euKi3ISuq9mJp7mYuoyB95hhKocH7EqlCv96NsB
1VTKT+2MZcqxuQw5wT2BvbsT2S4vlBwxpkpvq3jhEZ3UsflOvoF7tFvcCyEsJRNLwR3xIi5Bzqxe
sGFqaTpkbIBk62FtSNEI485oL2hTfekszqCud2/cZa0/KBRKUfTfLMVM7q8cvKE11Nx3U5+IAWwa
8EjIVmOHPueJ+qBAyorfbiUfhERY4Zmi2mwgHqlydzip/hC6Nic6HDZeHT6luIcZdqPju0vMqHNI
wTrmji6uHndMBvxoG/XyImPS/1lO+EZWP0BP/PpbYgIoIuKDG9nsgEmK/xprroKEARbdSQM8zZZT
b2VW7FafNmDVv1yEzp9WPvuw0zLsBg09PCPr/pSMCFimqFLbXkaWN04z4fDqAj2MpAVtIr5Dsqnd
ZmeET9fk895BVC4Tt8iKK9/XpjOJrukTW8PRej794Gq6oR+3VDQ2Bvs+h26x79ZBUrJl6X6NWxxV
uXqdUJGkJgu1xbiPfBnAeCMTdNgyXOWyT6qkYL9oRbkssqAmQ5QrMwqbrQ7uzSeOgIaGNGoigSDt
T4tLsBW9R6tLBHsk8DE1t8e3Uttrc1LU5owN2URsD81IUR4YRY9/i4XfymclTAsie8fptbOBdvGv
nUeLv5jTBL1GvgBGNPQ3n7n79D/kdKCN6qiOGIiGRvvNqVpv/I6kpXfqo+nCQsqu+NkpDbFmYoyD
OOuNg/lfajRYvdel3QEeZtufGw26QzoP4twWrmZXC+JCnah52OTOetazf5ALHn5cTjm6kmNadCNA
YZQLp9ODt5oiEAzTVWjXm611nvy72MIFr7Br34f1ffw9eLDE08ytQ8fMJAITmq7NfQRZv71B8+E0
EzepStj+UvS6T3Y7z/b/8/0M38cBF1Z1oB9Fq8MQKr6BOFMhLsMLWLwini4jbq4FUGX/3p4wN4GX
eL7xsWKMSSSXUsmnmfajQzSOsVs5+4STLY7mvIh/lR7t/rlji2LNqFcF4DG3m2OPDd6kqhkEF5/D
xORjxDlIGxKce14yCmbSpv7Lfy+U83GvqEHs0+ngrREFcseJFMTStuNVgbd/LPytb3bJwzqlVCSV
T+jJYUj4y3/iTcU1bw+b8ko4xm+Q0TPIpbTJz5ggh4AyJHJox1IJa+GxM7eWmSTnfuW/bc8E0dvv
Vft32KtIgvhmwH9HSh/zGWT4GW4GWdEHTIdGYpitOso6xzAFgNPAdydatZmujKmjTIldz5BmWz3O
ltPDuwojTmV1J23HTw4jVQ4NH6jQ9oiOYB9vTQjwLTE9jYkAu8Qly8nzEH5j8kMFQVpna7DxzrJl
og2Pj3sJHvosH9kGnuaPG6qI/Tld6d50hC/3Hu4gL7ByCyuGTmQLn2T2WRrMtYC10KSKs+d0ev7Y
2lbzZJ83Bt8NzwzTMQDaMoIrrG+yT/Q/Sf11q9WWcMsNCK8ZA9q3CVYT3U7K/AmcjvsrasEDXTd0
u53bnWB1kJB2VpN0qUO5lwYcKDtEcsR69Z4Foy13TyLYv0JzVn4StBEg3YvVviPSgEaG/CH/sR90
sRJUtdMV4hlepU2xr3H58boVlkESOoKq0kEpxa5whcz9HiwtURQr3a1qRDDxczP2UTceA5rxLthi
NAzE5t7SSPfKMYdENmXjZWiaJjA6RFIVyWdPTyscKKqhLZRznHbAXayIv9tD0VJBNEhj6hZLbOY3
7jlbwJ4qn1hz0zikWT8lHi4z0+u8vVRAFDutVr9eYF43G9PmJaxMG4nAo1Kj0Ebgr15KIemRfzmO
XWR7Dtcad1N2m7+HmMOWQnTuTP5m/tkPiP+JRaMdkU4inUEPAn40545Cpt6ERFX5Hw1+/Guj6EEO
5G32b/RDKCc8FEoJZv4i7c4kALx8QzpCc2PNrS9Ku2Usi3jiLGxeTN+vjWuSWcJzHa3mO2PrcpSQ
6Ko7Kc3i4Yj/4ppaZZTi9u8nIU5MmByPqqye3WBLPBHTDSjKcIqVjgHm3WdutjCdqrqeGaeLiiHB
TOyWlMB8mxl9P4TV5+iQoxWO9X/xLIQaVS3qnrVHI0p8T5rYhS8c2jgTYWZ2qAYftwBhCPk+Af3g
+y83ZcUNmjCwOm3FYmOAVT4bhL3bFnvOnPt5kCqqoOhT8I4mGk0ypguF5gXQwci1WEzqt1On7HA4
d8AYoc1Sk71FCJesWR3x4uYMkaJzKHHERd3YUEHkidrtVpi6q717dmJ6LN8NXbXkNjrnSlHj8cT7
7469Zjj53B//i7NW2PQqtaDOQeZLyDhwUubrTofLYLmhbgoZexgrXEhWrm0pDpHkUop5VSSxmP+2
uuP0U8tutugeB3m29YQY9he2weFT+IL4TUfkE1U9Dj9qjtbCTDJi/1giflQe2UfnNJ1h+w/CkRhf
xZlCY09k+jdv5ghXnPW12ZUY5OL7FaNbl4YiRNccBd+pLpMh8BH6HHS+QgB1nzg6SdifOzZ1QlAj
JpDrwvV1aTTjsU/+Fq4Z3ihWV4lzNIrbc7TuaFn1nRKtS5cSulj3ZeP03Z3Kv74ygeYunxibdHlI
1rA3vdXcW1EwEWFhdITPfeG35WrAGB1I3EiRrYW771ysZgGWZy1KWSOrWRrhJEGNLVFUTCCf+zoW
NgXGJnaSAmge8DPMcAhH3HdEF7T+J3Ml4uMxX5O2qK++tp4Jcup1OwMqzbvZLOoXf8b0INd5ZEYA
za+ntnjirAWBVowFvwszuTOtE0cUWRaWKHJBW3LtvAgq/mExdvaCVwMiwwY65dMTcNoHIj4e8K6m
zVMgGERer6Hu/uLvxMExse6o7sAzYxOhXV4EODWjwW3YsrhJd3UhQ6aEWxOgiNK+29IFvSF1/EtE
Nyvww1K1ySg5Hq0/mTeuZ3YnOXIXC18LTnRkyrhxmbz/q9C7HJQ2PhgBE6O9NLmCCXzhLDtFvuh2
9+Wxrbc4kASCIAkbFxbdYmpP0jL+0cS956GZU2j2vvMHKn/3G97UGUm+n2NVuvdQ8wYxibUzqVVp
DTpsuozGY9NGVtj+v0iR8rmpaucdL6QRby1ptU9TETYSkEaB8mN0x6ghqWWvL6mH3L9IoTEX4VKn
mg00VJVu2HpUC5HUuFs2oAiIBlCJPYDnJdRQEXwDp64RVn55Zf2MnC+7VgkcB2O/YL73nJB/xbqw
8mY64KyjrywgXzBr1h9Ej1VYV7zjnbt+pm7UueSEivnADKWI6Byq4P4Oocmtq159v+fYJ3xEg12Y
kA4tDmslHbGnmD94RV25n/yo+U36Eglj9QaCAxvFrF5Bq7LH8oovOvlSg2kfKVhBID5CCE2mN7k4
rd38iEw5IfFnuSxd6q4pHGBWX0BRPwuzX05SLU6QNIk/SnA/+5nVKilmbGkag7v/3ZkpXPD7/n+N
cKg8Rz57BcAU0JTAqezJiltud4mrbWNNgKFH7L14Na6VHCVFy+/ZcDGRg8s2TZsIdRG/6AcQXHgY
H9hXhrcDEEjeqky1sbgnC7ykbLuW+Nm+573dfWeAR1Ai7u+c6PCcFeR7+dFsrcytliYZXh6fMHUq
fGBegU8ss6JtY3sSIO01hfg6G/PoN3llGBu1dt/cjqolFQYTG4dnXbk4rptO8j72mXYHnNpHWmpY
0WaIYLYq9/ThY2hlxsPsP6SqSSMXYus1PKhDzJnayBrUHA8gLwarJ1ODWge6MmmYozhK+zzIe/Bp
TwQBsRc/pSoUxZ5iw+mqeFajxDqKJelw7Kw4bpP+hQZhW0hMJW0UO19Yw5OZP1cvds3ZGcyC2Q/f
prqGCvZ8NM0iIc5qbFUejNjnKkdGw4wzzCg2/xSJgoXn36l2HG3EJHrOoEhEihAPtaLpfDeS3LYQ
CvUrpOOg/mo30pdIp/L6+BzIWkKWw5BaDQqj4bv5xn6+01QkOc04hTM5kxj06aQExZD2VtWe+lo/
G/H7Tyy9vqEm3UiD4Wl4TbeF9yc1TU6vFDxAGMXi6YkpEZLMOmfvxibpzRmkD01D8RwHs0DZBIBR
y87qBhYpccouMYW/bfoNLqIE+Du8OLbG5WUhp1255avHg7ekBAGFOz7UahBYZ81ASU6TbGZVE5YV
mUffp7S5XeViKZ5iBDEDAHkzoEDbSf1pU6Xb2DYKAqbwfdiu1rG5KaqLbHm3eJ0SbrXluyeUxXJa
zg0nJ4J/TbTzBqQc7dm4rTA4QBLl0CwvFP3Dd9YWVc9Cpgds6cXfPH/iuOSNqWiIuy51ZNuUOEpH
LBCY14oEYZATt1lP0vtCqoW1VBDOIY89D0XbBHSBjAI86b/N/anLorCS69j6bmUXzd8fibXVUvaN
vmOWpaexewK3eb8GdnV6KfgAFIsrJxKIWYt+V+XodQCmKrPvM5BgGZSJgQ1z3GxVQIuizrPErRfE
Ivey1KYtFDHVrwD7lq9BJsQP9UnYSK8kBqFCvmldsc8Ql3q/VmLz+9dM+5QYhuy4G4DEBc4V/k7I
G3T7B/sEMML8e8rqvI8AMoCX8jF96stei5mDJRgP/jjSX65sz0uOBRDBcTt7DLwQ2W+rtzH1BIdg
l9FkewHe4/P6PNwBvncXIZnkjb6mdB9Qb+uirN3Or4WdQjg+4qWRg7A3XIXvwtXwnrOhWVIDUqAP
C29urJd4pvG8G/FuEThrXAJ8fYaCjV4r9s0E9FclX6Op8Ba/l5XrYMWcv2O0In/mP04WXodnaU9a
TBg3x3c8iEqY/KDqdQdtR4gYPXJPt1KjPaeBnS+cRTmMtzmx3dBAZii3OAM7Kbm/qYmAmXwtVKRD
9KuxEB+TGMRCGAUnNiyrh+pEZt3J7UDqKse0pDrQss905kUlO1yo3/O43BSfASV16Pc4a5NA7OUN
0QnGsf0JNbqB9MvLIJzEIks0HFuQIs27BV13gYbqIs4PiVPjVS36F9FiWZFFbXGmJgQHrwbuYSyu
O0Bms6NklndVVg1zeIk9+FjhdS9/sanhkW63Jh3e+eR3IkIhg+pDe6Wm9wtKYeH2ylDSbMhClECh
lxLP7hXu7Mrs2kOUPmmPqynuKshVSL1Wv28eL/AcKbbcxbVGK17gEM6ysDOSvtUJmD9CIoNWAACK
ysWBcDqxDs1DjXUXlkrEgjTEbDw52t6MxXwsdD3wIuUNS032T624S6/fjng3mhBcZOT1b5rHwKHc
5DcEmXhkQUjamKe6oZmaX4rRetjC2pCBnrqV/dFAcePlr/Bug1MlRgJhncJ5O0P/WnS+Gu3wjcpn
+GskBEmjFMtNoFm5WkgaulRlAbD3AqYe0GqJFWZjykHb1VL8LV4tpAtbrpJrcEd3xcxM3+83GWq+
GyR748hW7LhA5wY5S/d7ONwIPzeuJi12YGvG61HyvAJEm471i45fyEH6kc9hZWkrO5KNbHUEC9N8
MYUJeLerI/7lzQrqlIp2xX/i/sXsclkM+MJ8htGmhMA6+oNCRMvT+1HkcHG/5WOHj+WIBKPnC5tl
y6/KlAsee91tj/Di8yWR7kePxMgGWtfUzFmuA3Dr+4TxTBxPwtbj6zWYLYpxTHFM7OBipB6IEuGq
sCWVaYySCmxDC1dJbt4c13tOKXzwdOxev0TyaPRYPjW3uUqGQUpCnUG+u7TwCQtSjKp2WDy2O+RA
4TisUAcf0GK99hNEatCZSl9NSXNtHUebg8edzoQxRXVaS32xXoO75J0dfVCEpkXI0fyuzi9Ih5t6
lDteLSMsSz7b0aRUolL6+IuR56LVvzByHSz99w1vZtKw6YvsoaFI7O52Ad3ygoEkjp4OXvDzS7AH
0ECo14rcxvkxMorYlpPw/uJG7i6Ea7hgm67Y+SBTZi4CFxVCu6kURuSp9beYP4gLSJUKbY7M1ZBV
UMsvOWTwFCg0i4OVyyQK5WSTXvb2t1Nq/DKj1OAUqeYPGzcJolS7mum74Vxces5cEJgqyxF32RNu
3g2mC02iv44c2T/BScl8AUREe8Hg6F0OzhmpO/ROjrlILeARwBbtu56SDmPCNPAhFrBo1Wv6TFFD
I6ags7xvwYxQs0ZTOPJ5n89lB53KW6lONHjRyGPR/W0ztEB9rbpf/NTqx6uJspwOEsFj3mz47mX4
s0Y+XptdVJJUG64m6dKBAxTU+Z6sIeaiOXuxrAF+kqPeieumQdKWL6dRSweOEIH2ArOAkbWNVISk
F5+hodoVDjpp8T1RaYwKcdJqdRQE1vjMpOXvA3bBQbtB60dYR8fWu1e+OJOKfr+nHJcx+3X/MPvc
nEh4AwLF+Z3j3kIl5Q8u4I/mi1Rkxe1mBE03jgSFSbcw6nButO1rq9nyBhEQQ8vju+Zh95nF0gLk
igno9AUoHxP/e6iK9WfOpAF8CacyjVBpHavZQSB5N9K7Qz5NNJ4/oJW4/AxH0e0WfJmRPh0NnfFQ
XTkI8lh+qOYODdXhYA3hWvhCM+Ld0P/iEFzN8Ul69KdNQiUOe4RxlGs9seEiSIj9jhjvzzH3LgOV
Ka7dcjxvPY5/lLYSca/Cx1CDdkbY6Pyuf2Q8kDRP0fygssep1gofMU87WoKeVFs/zPScwjB6BF+G
ROWzjKOVoe6LkAsrODnLZcbu3DhAeg1Y0xfGmGGVOeKBD6IanHuEQS8MZG1MOjDio1ownHKUykF3
jgb9mN3PKJsjUxeupB3PU5tfQgHOzq85LBq2ODKAGTtCInKPRXljGeATMaKxezBVmvdosHJa6ZLF
GtXOW9DrOQDPgk79XI8F3WRle1wyhnRGejw21RXZGlcn5AEMLkwh3IfykF26O+fA83WC81gMlXQo
sMWSf415voV2G8xM1qGFEGLLuGFKXgTYeppxL2Uz+Ps4zyvFwxKX3WK6dEfkuB4uxecRfOA9pMt2
XVWs7MudG5gzmwf0SgzU8R9o4u87n9RzB1rA8JHo0vtyEaI5cCNMczjWdZB0lKhknI4mHFHWcfNe
MVaQzP2vfHp9/zpLdcHqsWVRW7dGNzZYSANntBryoMQBV0kAthjg1NX8aAFOhnRtAdcT0hu1ZPLm
/6UIBCZQMRKLom7GZafUaDPhpp+X2AL9C2KjBY6Q3rWJTUz6iy9G/wA/BOt8JWLEtB2iN0ZKOP55
NaiV4QtBqRF0OsC6tF3bGpD+fvQdPn/ogySzsJBYPttgPIm26EX8mqaqzJCWzntYsqYOXyCdzQ8R
uDylGKl75+F7q75JtS2P9zWiK7s8WlvKENrrmMn+jamMzcJC2oNizJB5q/sVM0ebmE7TJSZOhzqz
bLQ7G5aEOP4bHy7nM2zm6+yPdXuhhNa8OvNiG4TiqMinSFcG2gCKlSvHe3j9kmQFmf/315jSFpso
V1XZbQBbFP2Q2IHryaED8/TS67hZAxBLTO6POH0IhyVMKQkNibqxyi+6x1B9nPwlDlWteg4YaaaO
brf+fwEXEcpSy+wC2b6f/i4W2BF7hbzI8HVve189inyptvzqDirDbXXE4ldHSaFnM9qPjbDjxyTU
e+/TPRFDEgXnKQ6ZwXIb5i22hQzFNeSuGANla1ZRJx7bXS8SbkIq5dP14XnGnaU/A5Jv5olzCai7
55l93RNltQtRwNnGZujlATeD2JxY5a7sIy0nTuLHOI2SGjKI9hPK2nt3BC6cJgb0vWIgyYkh1jEA
meGyKejLkvNOFZU+1FzCKiJmba5L/oFlT6SwrlOuZ6m7G5O2un6P/Ck6GspE+sS039efcxZh9ctH
fqPJ84seVe1ljz+ocjHuT7kyLTJ2kkRPor84eBsfQaPUBJBH+TW1sy6E7BUFnI4zoomK8tBZuhNU
TgYQ911GoypB3mLXMOj979tWUlT7mPKno5oYi5MhEzdKVoyAu2rJl7eK0N20Vhsx3is9AUQAzmDA
wFfu3awzE7ESwLHLepKeHywTl/bsJG+3cSfqe0Z3+Obrsxy0r3sgk15OjwhaguzmdU8AYbVfzvQf
qvtkA3KHsRWoT1tQlMqj4pcT1RuNW/7iwTLBXqWl3d34Bm0rmH4r5wKwkGzdoRj2UthFO6na71Ss
XwZkKt8ubnytltInyGfM0RTWIGSuCU9+BzuEf5YYTPUEAc8m7cCOUXNMh85L6QwliYWx953yTqRr
kxZZv7KB4q0LMwHzuE+9crb+Y6i9jVe0Hi/zs8twLx7+NgQBANxMRWIKYAPwIQW7L+2lKayERFxB
OP3TapZj0WxA+tmMzlHE9UXz8xKSqIOy1KgYUBBkjL9Mv6gorRk90znusrREDZuByvhcB69diqIc
yq6WcdU+o88Kkx2r2uD+P+6xk6sGinZhM0voHoyG8t46AhJ2R+leL0ff0JJPK45Mjr70YBX+FOWe
Yw59nU7rsLAKn+AofuI8PGS665qXCKWrkNrdHUaJMYkiZnqtdjB80ths7+bxXr8pRporUb8ewPV7
K2CWo/vjUfk5U+JrUYpMb48bIAtmzczAN3Q6vXD2WdHu0VDLL6gWY+XeAQVnEr69Uz82S9Ic5WhO
9N8QrbS0q8XFmPBOUhrlDkhCa0mkUEuJhDDHmziTYHM5rlelW5ajZoU0pZjZca2ffIEuHtC/dmaZ
mk+qW7ONdeRTaJLMe8D0LTOwioBUd366taBbOL+aynhrADFVG/0kZ7aD9HwK68mYsl4i54eTduUb
O8JdYMCmQIWEn015k44qriBvLyjcoERbsk/Khix70Kg1H5L4lpaWszCaVKF3kAPSY/197UKTAzYd
8BXf1zRygM09J2Bp2XuOxhZwx0aPr+sxnmFJAFgAji1AXWXDdP6r/adzY2AjUP6Fdeg2G6kYdgFD
4WKOVa2A0yoi3hfsPLDpvr7VMflekWbORxhBbsMtVLsfyULv8ZghFU711I3ZIvft+A4EEP0PQwrv
yY+BfP8TycTB/B/sPVua4uOaueSaalJcoxmBYi+xcVeoLz3IEWllH3RUf/VvXDG1rRFIvSjhf4pt
8GWfxqE16e5ttJCw1TNmBHwxLq6ct5rCDeGwfWERc7qV0uIyFJZH8yHOlPcNGRoenWrKS/zzcMod
8WTxymvIVP+2QzX4WJExyRK8pR9UOSnSW/QoK6YPVaUn4svl6sP0JRFoCKiUYw8br04DmYRoLBqZ
duFlObuDvDNNCo4Xz1AZWR8zZBSvDK305rcYO8twglm+m9Dys8hYNMze9P43Ivh0dkJf2B3wxIer
mZYblHLl9RR+If8WSmXn5FHUEHi8M9dflpE3y0jbBryrOs3pd4B449DaX3gTXcWSQN+rr71yzpRa
75Bcebxx7/Km7uNsCTLLUN2XhFfgEPSBdyPOnwTb6W9vDSgFwFD0T90bee4kuBqnGqqlgGIMuaFw
bnJ/qcOSkp22NU4CJyt72levf6wwaw4eDTofi+CqGiQGdyjHuGh85960JlNRFNHryZiJGE76auTe
1/AFFMA1FraDLb+bl50jUjbzEPB1WLtH7LZKU0nkhXqqvD5inCTo4OWDNJO6bsHqBLKxtHtr3z8O
vsK3t8IaxAOgUXGdaYzfyW0ENcHcl/c6sibQ2g6Yu+2v0xYpiQstirGi+GUPS02uawewU7cADDGQ
QRescUJdlIIkQlISAlEWd1ZO1Q72aJoTZCyeMLkeB+c9+13jxX3pWpYETFclpSs7jhBl5tFBhs8/
DZbjJbfoqOItFRpxv6vU6q0XA7sNY5XBJCuJVDbr1h4cSI4wcwyalIADop1rvfkJlU3UCqqfPFx5
sM3RS/ThrY2smwDK6G3wXiqA1CDwNdvvAzh2cwjQb2JnLtI1GwKX+68fmG4kipll68wWK02h1QfB
peeVcoQIEVa8Dq8YQ+CR7/OKjn+W+A7TuOstbpmofR1pZPagpNgk4qHyxsdSVGiOED6MBLK7BIU+
JJyX1iRFwn8Cet1zNe9hmGI4YfMJ10a9pc7K7MUrkVrQhXzazYf3zSRsGmqsIb0A7MTXbdU9feVb
zUVtXDwUduxIFDvxIa9ZCmCjFb1DLjAmkLRueQOKPCTSzXWUamBOxKpJTjSD3w72P5Z/OU57fQgW
W8wDaLUEcQaun/1DNwJkPu4mljUpb0D4oYNHczeIk//XmwYf4XvbkaZESk4T56bAw+/Wvu0GsI8M
ArChnKyuwlRkmLpn/S2BhWVJZkKdeB/0lk8YaxLzn6Q/Cp/1uqFzvnDJ20j0RtFJwHkaK/lgxDt1
lrq1Cv4VCTJ9udVb/IIBIopbmKluS2xFMEqzCehBJTl6RiLghf7uW9vVMUKiDC6DwNJCY1tppU2U
LW1TB+IMl3DgE9IYb+SDpL+brnOo063oDP1tY7/nTyNYdI9hltUOsTeI8N76ERDssVhyCqUFen7A
uEVJVCv40ODX1qWDo2bmoYmWHZB+BI55fMH/tHli5XFl4jyn9hsVX3XPBO900lTRiGBoZ0g0LZEC
BbhRzpB/Qbfma8HeJ94r8OfqgPwktif4WSa64hVhUmaM7XWysij/RbJlkob5S4DArNWvWhlfAtLN
5Ec+Kg2/I5IGDV5KvlzEPdSi1PbJifcnD0+QYPxCkGyZ6DbdUEgXOVrG1bERAB0hB1sut0J2CQTW
05i8bLJWcXoHhiQ2cNNQ97I6agp6bJ0uQJ7YNr/ZxNDSyrsV/YRIs8EOFct6sxKo1DJ5t3USMSMm
u9YDsXwOV1PKitm1GqLD6iz3xg53EfiuawMuRhibqudYEpzkh8Fq2VOZGcRDQ/iBhM8KVFmNerzm
2na5jZBTE+oYwJWorBJFKCxo3jrAJrnesOmRQDLB/+5os4qTNgCgLoRf7JBtBpdpkFf79sbutKXR
sv2pLYznr+fhG+Ofq0EWAZC9V2Cxl3+8UZKv/GI9e0doud76NIqgaRtccPFhnyjpggKbpACfbyfQ
Ic2pAfcox7i8bVnX4ax1KmTJEgK7DFiYCufliqJA2DEt0zKP796KH84IhNDwQqIyB8D9M5qxRZKN
1irNHAq0PlLGQr84dHYIGvD7NnG0tvYBkfPLW2vbrbNZ7VKYy1kG+CDYobcZbGxQb+cpybZwDZAk
+/WXJa6RMFLUUk6nNU879i33NVaY8tsRb1oKDXMth0oKIIV0/g6XxZ1J9S2ZDqpbNjQEPWJe/lV/
ZqUYEeS69dOq/NbhwJpv9mAqX82H/axrc7IXLlv4bfcwijDgIhfvGMVtrvGvjwbW2+5mjPB6eFXD
/qGf0efqAp46YoxXT/crMpzwV1I3nBGEhTv7vjUdxnsA56vjST5NpuLxS8XVvrOLA+kzfjPn3sWu
IjiEPX32h9uyREgQQd2jjezYABNyqGpNVtsLYB9Lwt7qDFkHvuElfRwBJIX5+hRfF8tu4VEkQQ7m
/98fIy2WK6OBSOscxChOcGA+cjaIA5CajiTGTa71IN0sSuKMLCSBHrLxNEtWHTXSbaU8+VqNoJET
wCOO7DCM9lrcTnDSpfYgLgdT3gZZF58T82d5IGuRVi+YbKVVFEmbEqC13NosLfXxyF3Kn+SGPsK+
+rUoGTv+POero17I+fz0BxkQJCvqX9n70H93i9Xsv25EsWzoW+vIpyx+SG0XM+nk78xof4Ctb1pP
ZfvOWqA5Q+MEU4ARP2/lHPkeaKlWyKumpT/cG8v3i5DabKrywQ3652yCsDUAeArdHMZgQRAaMSAV
MILkaGjshtm4yQz62lKQ8fQunB/286lnL+ETOTlhaKiV33q7SUzNZp3PDdj/jlS19pWgcae5eDOD
EUxyAtlABmpRHYpfY2PwYRXeEeXVPiDjkBF781vAI5lO4Jyjn8siciZ9JAvGZHuaIsZ9qBIFKhsr
P4oAvA1/ehaqTO1mFlKFpDBQlhCUevEDzr20uZXnSCXO3o4cY0ANiE5Pum8yUKIjqtYStzHCBXfw
L1OCMAtYEARz23Dg/aPtqVWqg3NndQa4lH1yzXQlb2fQyxEuy6wHZ0iOOCEEOU9ddKkrsL70RNyz
U2vimHHqez4xdLV1HrNoeTYPB74GNul4XVseFXCU0RQkjdPrj8sFihO7VVBdnq/+6a07yn3yY1VF
UyAWOWItzcbNrFPhfaDGL3gJtkrY+TlGVPGoqCOmrwl9URF0h9Q2qW56wWMv/kwZ1WzAbS5jn1UE
iEZ8vU5JKxg7B+Q76mhYe7UkCp3nV4Kkf9FKyCdEfcW+pQ9WK9p1IchLBkXo9Lj9f8hYwhingT86
O6z/1qyBut6HPXq2OTrJu6Alj+WWsRrNsTLy7ZXEash8uCTTOQRmutYoigFpHR3fWkUw2gp4dqEn
/lPjykqOq0zSgqegrCJY1OqN7kVAH/MDefKxS74E+ixz7Xt6CRnigYpQ9Ou6qM+p7bjXXVyqNkh0
IuDin/XsnfeGng54Tme3D+xOJ8IZ+NVLEW1ETOIFR7c9rfMhfHJWRGbkrZCbgZoHfSlb+eZUDyxX
aPadFFxkkw4uzMsx05xyzSlIHTxXpbL+fnpST2qG85UXi9jvFbIkm3YDhZ9wjSctRg7Tl8ivMLKJ
caWaQzF5x8EEqSnZbYEK2dOmsaK9SHtDBv7F6hOoWIPrN8IUZRec4e1mzyOi4rEuPIycNou6jHw/
azt8Ozn+jtRjJFYMYUXmiwBWoHZP20CEujSb7aBsLTvPT6FH8/CHyw98n7nywLO3VMjZVLsqfwhT
y1ufxUDPZLCAtBt37/BWeexw6OrAb6bF0uMaumDVp+s4DxXr430y02qvtqGvdNmOkZu3VB52Jw21
ij95lV47nLCm+o58HgAjFnX/cg2DhuSiZSxL/hI9H5eOcO4HsaIVoQxZrdrU9HOmPjz7TFxNH6n3
Hnw82WGJR+MS4m9+0+oA8Wk+LjoJr2BXMnua2g7Z+Lf+OgD86Vq3tA3Yf0VVCFiuGEBrZiLfS/s9
T4QX4c3FERS9vU6J2NBi9yu4mK0b8GIoBsg69+Tex/r7IGmN1Gsz+xBE7Tw5ywP+1aaXXKqCaC7y
LuOHSyICkMyLem9bthTr5YvF+7ImqPSn8k4Rubcc2mwz8LeWBA/In7X8G9oXPehWcFqGnhPz5+Xt
lFu+f1tWKzfLU6Fnio1NLEX/F/RckEA53tZAJWAIm72sbOhsvll2WCzej/P51HPbKAH6ciZcrgjW
GkkvzxvIF+xC+gymL1cF5hdk3ZslAe2CospS7I3o4x79knGGiJv3u1wxrlybG3naCmhtfWpEk/gG
HF7VBL+NdW5AMsEHxgVDViA8TTZ/HpsH3bIbKMLABjWky05znvnDrD1zOHDMlR6PntQe23Gn6B0a
D+U86VjT9O5xTHEZLK8xwCyyafihuRBaUD8BKozYo03PyQU3Qg5m4P8+6yvotC8yU/hKmNKVQJbE
bWqDAZOIjLr8JAMoSUjCGD/wx1R+OWOPIm5PcSiAVOq8nXzQhnSoaW68RrjpbC1xQ4kf6/p88QGs
UW7emdQbIYCgEWT1ylH56ONsINRcE/cmZnHb7uxGneLxWHHB5P/OldB3udRzh5ZJYizcr24sOA1+
csjXNCQCIiD74ZAxDlrKMbgeW4Bg0pVx27ZcaTzIifA49HqnKxmsYRguzEjfeepSFibv/l+NRzRO
xc/e6B4AcH5HhlIGR99eGzktvQbmCSmXiq4vEYyMaHdf0dsXjiswQdCeLE2uk0jYbvAlSvraokaJ
3Lo2f3GDwKgvlyivpDogJQOvh3W0SrcI9mNhZTS4xWp/At+rPRX/D8toaryPHodbpMciajtK63fm
cMvT1A6QnHPFZ6gsm69DCxHqzR88DowD3T+NldoftmdDNXFacHCmaZpfBDeZt5iBrTvIb4obfAXD
ggoKhzuGh9ypu+9tdkyESoMEBEksGrmiJkhG8aDhQrMpXsk5m+cDWEV9wfWA9EqX7YOpABOaLvwG
b/p6yGvumBHyg8rK/Gchg/9VvyluRES4D2uhNx6D9hd65I/SEGQnq6/khbB/JwVmJCwMH176C8qD
Ur/6FDTLuT+piAR9Hxq0jhkfFTYDNV//Co6ZdISy9iJ7Cjo0GyxzOT/8+kShWquq7YwGK9QTloO0
Sqfi5unWiNLir5XRP5gF/f7H4P39hEXaVFxAZlkzjEHTSIqzBnpCskL0KNKZDV1V+gr0Biy5PamA
0Wd0xvmwco+Vya1V+3oTfHBOw1DGOdRPH2YEDpzgwLAClKV/h21R7iaKVhoCR3miAZY9Sl1QiCpQ
obRKcbUfqrfHakXxx1uv93xGaE/8us68qvVKtACbkhqzcVhql7BQK442BPH6lxrLVCtAUZVxR2eS
WT1o/PThKwSIUXPiNgcRFa0b1EvNVs4BtS8CzjjXElwinvOmDxemk7Rrq5BSz2MYh6v/A2WzckWp
gdu7I9GRLIPLB3Auklnb5MYux3qgqlsD3DEm5ztnTdm5LcEmCulplptz4xdUq6eNucOUJ/r46Xd+
ufyYNN2o1ryTVnw6cMkG4v+KqNzbYKbqteCAUWAdoaycRzRwygQIJHuETXWbTgXnyHwTm5dj1uhY
Savr6B6ZKwwUrNvclK8n3DkcR+0gUA/25ZUXBWznAgdC5nvKxeBVfkO7ehU40NMqNg2qAD+Uvc4X
t62e8lMoZEMM2JfwqSBBlVMe8wkP23Cwi9KrCZ8wB94znGqcbju03+mJJThiBe4lBfpphpUrVkJk
wZVnM8Anz+On56Vl2CeScMlHKmyp8XQ/A2+lPjZgzIMIfSPwK5+kTPoY2D5rPznda56TIamcJU2y
NdNOWaILN3S6UuGwn1KNRPr+8NI/orD0tOzMx7GPDCfCvbriPxxRYr5AKX7lM1gzawnGhSyBx0Re
3h8TMqpKLZZFpXHA/vYnVJtx//EgjMaU6ipj1aXsa60IxoPCnUyWfG/M1LbzjxM3YCp4ORi9mM8L
N6vk019c7NDSFBds4DRsPBEfUMzSM+FeRqdyv7Q4xFVvug7uAFJQclibsuuGVGKGulICECI50aJ9
7vfoGY9x+s7Quli1aPeZdbh80KlGWbmhVwXQDeRNNa4d7wEFiQbZDdOAuf2p4k2kAjxWvqEePlLu
crs5y3ZBdahVr8OBtJ1pqGFkJZFf5hzBMVDPyNPpLSI6cTYsjgAJPy2l1nB/NzqJ8C0+oClciYl3
ZfIrttEFLiQ00gn+a8DA7VYcA0j+D/d9BJom+zaR6Neg3g8UUAZYrPpoOKgZ/LnEYTpBjoEaVCf5
qR1quRiW4mL+k9gj2CtkrSWUqhUj6iwRMaVQbb7HZ5u2rrf5ESjx7BxeDV337jytn3fxAOaefhSr
rqB5+ZCHpKfK060Bg72z4Ezbfz7wTvp3xMS0FTFt88NrrGMECBKhrV52hDoNAvxb7UD6Qd2A4qbx
gx6wue8l54qYigZFkUIYRtt6YrXs3vE+/AGpF13dcQhsXaFi7MZUC3T9dcpxRhAmL2B8Jg99B/2S
MQphwTyf4lI/60YJ3atzGVDIX0tP3DNHforb/q47gXhfYphLbido8RbGO6Jjhwx6eLulXlSXh/Iz
m4IcunoeSc8NaBsioS2kE1vm0399CUbIYXriBT+ekKB1i3KchVzRrIK1kjK9LmhYlec1vbnXNvlo
sNPFtHgZV0m2dAVhPU4BtR2FZOOTyEd4/NFDFD/D/7YP2YwzJz0ZJ97cOzAB2ADrpqPynNcOy1/Z
ftKUIHQ4mgOKbFMnsuFRolhL+H58bMthce/q+IhTvw0++UiX7CiHiDqVv/UFLue3DzZ84Bne50Cf
uxn7nofwceEf40+8lC221auFs2ilD6VRZ5at7ONOi8w807r3Sj3asxHOZ1FMZLW7G7hgdLdnO6w7
7vosEkqbIFsTaP+zvfL4k9ls/HYxCRTFizMiXnVckdrCle0ZdshEb9JeoUkvIy3SNfbI/UV7zvE6
FSbtWOb3Ut6w8n5bo8bJa6IFrb3RkUxGQvs57YM2ngMAquHMAThrffL3AvDRT2oYp0zxPoU2O7sW
foIQbOYdpLa29OD4GvlCiRVgyR7WHlhKtiUkRTaNFM0b69VsIoobzDbY2ztpqSmIUsJwUY5oFc0j
U98zMf9/hxF36RYgBHyYhJ2SG67b1XK8TEYLwE6Pa4WrTwmWmciTA7LcEYgQ6hZyikB3s04sGOwO
dWeaxodvY2/MCUvqFa+BZCrKgxk2iTwZJOdr3z8sKm6rW3M73fReXFFhYUUdsCVDdXKLibetOsXI
9H6LFaR0kTwSUGof/Gu0yz7a9xLiXQMrl5inVWu0h7MoZbr3G23P9P4g5t2+zsCogEzfPYuj54Ly
VlIpVcOwoKDDBFsNvaEI0py8RTvaS1mXMKQt6CCU2eedDnTkiCAz0WPlBjk1kSHy/SaU0zdeOWRE
Y6ERnJCuTSLnCrc51VAeOCfPH4LrSBSRF/DpI1aMFV/2jNxnIBPNH1Pk2HIHUzZry3XzpHUDyoNg
RI1NYZI9uRoI0l8zA+0Z186FaMs6fjDwieZkNlDjzyk0ZUXnCr7vCLV8tmen+xF2R+4JMJvvU74F
E3atV0WVJ881tmrqzu5WD4B+zNGH8HaJrQrNuc0wppd7bnLUWazOAtJkuGl1CmRmsn95gqjPDtFw
o1+SfZENb7UWiOE12nh402omtHkR5Ud0vzsPGgOQqZzTdVEAh56mQRKYxefCkrAPrPfXQJ6nZAld
+Yev25KyfdOXN/+BStlyDZ5i5sGGX59PwJZnNFhoQH0nn42Gg+/l7BrraBeeIwqb3sGtCDRFQyfX
2QaDufhkdyt2h3OoAoZ72gs8xhDeki3s28A+TL2kGBwH09y3ZtDVEDuVHnKyN82XNaqnBMC2x2jf
g51UDRIZlsUXcYW53y+oR8m9SB0YTgiwrQY9LASkN+Dg2/ZjJQkz01+gJ53s5OqajnFH2Ti1tlMu
Fy9gsV6QOcXQMdxRP5tuO+kutdK1R6UXuT2MobOoCvb6qJGtL1mUmw/irp0oP5J4/4THsuEvEZyD
W1SSbSYi4RY6uFZp8r85UrnViWG0qh6mZLsa4UmBUwUJD5MJR15jXWr1ZPzKMpwQl4rkfLx0Ii8L
OE5/4bkDiz0336z1fR1a/Tx45SNHLaGURzZU5mLatvdZwe0dGmwBLQ7y1NB7N3QuK6ENfK2K8EWT
Rb/CyYecLjsiyM+lSGFYRcvrlWSODKZFchyJPmrO8O+Eti17hibUuuKD5FtZh5ITvpNeOQxeAHKE
urWWi4Aq5S7j4cvlYtSAwkTei4d8x2hui2pe8RVJoavGD9jmZnbKpxkGrCV7Nn6PnD7vM7cX5olb
p8+gQ44CCStJm5jj2sBKCR69lH+w3C4qFGyUcijGRUwdhX94i62DJ2/nkW9lkUhUybB1cWKT9Nvb
k5z3SThBQTPRLCxNYtWXoJX6UMYWlNGg3HKV9C04UwO1qLKWByJHKb+Z2VYIVoIasQuEjpj0KJC2
d7FrwgHCY3oqD+Hkl9khZz6/0cRKR9hSv2/BwaWHruH3MM7Rz6kSPj7yFWhurCsBmrderceOPdSW
4PvTtI1eXoyykQDDZGD6OKizQw4XMhzfF8AN7ynloLXMuYiImk9CnLy1KOKh+En0fTGPy4MkiSdB
hjCZIkeJcqcEFb2gZAW68V+tmieWpVZ6k13YtW9LjHT19HwRqU79/LImNtHXKN4Rb4zzOUPpg4W5
GUC6qjyQ6/k5WzQJZdRY7uJxE2WqzdmNHNkuAZErVo/AwBktLneIfTlCHliJuE+KAETylCOdLnEc
X9fZ0MVrBMiEeVwoCi1hIqLLUE3ve4xMIGRBQkBfkSqIXwMu3QRT1EPdoy+P2oPYrgFBjPBxC2bM
WjZgWL/EodRKrZK6az3wNfzBvMzS+CNvuGS6q+i3yHhwBZke5CF3hqzpyTXrst8jY5M87aNWZCdM
wVjDKUS9YtwqNBU8qSmHuMEzOQnPthmz1TOHlJo08ybajB6GGvaiBLSt8ZOpmZIpf8+NilHG104E
FO/2Se15vEdmrP9GsJhE/BvUsEQNcpWjS94dfIJ0vfCYKRdStbenhj0SqIDrHW6WA9Qynd+nz0jd
Bm9NwHPNmUHmDUlaI3tvnsvUE5QPDF4Ou6mYyc/uukOu/qfbz8YK4gYFYy2PbDpFrwZ3OmwQhaml
JiuKFWkUfzjzOP8qPofw6lkXWEmoQeDgGeLsluhfFyLfeySKxlMg/IzDfLykxhTUSiDNGkRl++5v
iXR2Fd3eWIDde2cLw6peDTco0Dt7tV5aWmGUpyv+9hiclgbqWjfSHlK6rSKNDrE3XoLaQyXak/NX
dXdqCBzm0QgOqZe4+4y3rXrnG+ougZ9xv3l/VE4BGaeTPrBvo2y+zvXR81EpWGYe0Sj3Nvdvuf+9
JLTAsh7C3MmX8FQ2LdjzIkC/x9CBjPLQy0EHwF1KPjwYab/HeQNo51hBy4dlPDkwWFtDruQsKIte
y2eWhiuBaLyM2sDv7LcV6ny0mmkOMzIRSOEYU867wds9aqEEmPgkubFAJ7c+rMxNaJOO6EtUojdd
LuMab0E651TPsUkFjSCmUgCvD6p/kQ2SJADy3Z2K7pem1bCr9NIH9dloVTqF7ew+7b8sG7EW31tl
0LR+tLKGdL23szrBq11k6gX2Ki3ioHYFpskgvUX268Sz2TQ0jydyoQMUn6rKa/m8ddNocCZifPHq
cRika17onnMPfSE5gDU4Zo1V4Bg587lEmUPkQ7cQDziFa/HBpBLm75SzbVs0OI+/pkkKM/e5ZGKC
9zIr2N/196ocC/XNN/hFCKZH67VRoQvVrML9DBCClCpb5mnzdzNsWjQkvxcUG8eLVtlD6cvfwC16
+Zl431fF3gDzSOwu8OqE0j46WuINQP7p5rvk5aA8sDc/bQlILlWbXNlmtoklxX/6r9OCnJxiVOIE
TKFYrgG3U8GJSz1ykFwcHsgTPJb4dhbKx/Lizs5W5KYGsCX7aVbx51rddmp+RvwujqSWbdEzYEZ1
C8zhzPlSnoaYIkmYPiWkjCChWJPYDiXgzh5EEFWpt+GeF9iGsaAUz4aYfIwnSFuQ1Jbx/INkZw1J
i2CsYh/R8YsF12oecKUSqfb+oFFWRjfUI6NzcDnZZ5CdNmhqcDDO6tPFDa2jtBuKno8nY8CDLIMH
V0IQIl7cgnRtiBFFYuQB1tQ3xRCZhGmGitdWNqSAJvBY/XPnbfw+2e+5an63fh3OuWIPQaU0ImGt
MU2GloEXyxzO1fKWA20PNgRsx//nyUa7bvbskDh5DWt4VncDai0lhSkG++zDMYf+UHNDJqKc1ouG
KOStIIJDkPq8d4Wdyx5xFniVhC7oysCJ+1IPYQLC1BQpXQu4Nh+7JiQhDz4NpbsX79anvk+imhXj
O0Tc4PA4bKLQIGawlo54AN66PuNAEZLBkDmfMw+PE3ixd1HSwN60vMV3qkdtKvym+T4c340z0Bif
ml4zyH2flQ6OA8NEr73gzxAP1bko+H0SYnPy6/9uqQVfKvMwowLMlEbQ/7CnJzLXJt18xuc/yYEs
IyKZp67dhiIqUbG+ZBRALynf1kLqlB5oyO5gIiybVztYQS/kBzdkP3Bqi2X9ntbPWdHFmgsoAlqa
dWZq0qpHi5f0LxXqbXi9yybw07d4ti4k278VSIbnrmMZ0MXQGmYL2G+Sr+H0hfjBwBoewmTJAtKn
sphMCJDZd/WtLEa00hegK0FBnvbAkK3ylaHG9aI6/ilZyAre/dft6+ruZSfzk1UdHWP+ZqsPjVJl
+VpD3TiszYkkxx9qbElI5IfZdcIWgX/k2BpRLCmA9aetmR0nF/lXo0AR8gUXa2r3EiYMrv1jNLqe
KQWJU3dI/RdSERFjf2AQk6L4/fwObP3O0vuJ0rSDI7/QFq5/hC4HzlpGE3xDbh+rXWXVrFgAOGtn
MRmPpML1I3z2pLIPgJX6+/w996mFoBQzabYSKE+gDiOrMQ+McAG80c13UkaKtT/qG7yrpWJUZ4lo
593OriMV0Hg4whj/S213KWX6CDr+Y/20x5/5z9RXRcYRi5O+uozykIDk6uMH4k7C+qYlxP0wybvt
3XuhXp2n0IMqbQqiXkO6yZeIHolAMWhS6vIVMuos6ZKxlJ37nvfIeOl3RessUYHTFHnv7HubF/9Q
jjEEj1tpqgsOuAHY3VpbBUJZ7fsBsAVrs486U3MZ+FHWg8obyVg7smbfEav1dzq3/9lRncuzDDQi
TDw2vyzpmQ+x7Z01xPA0aId9IriloO9wCiPAyrVPDNzK5CMw89LSBjrihjw1tKw+RbW6SyCr0aw6
ocQkkGsQakPCs4egGpJwYPAI7dhu2WOYVAwRTFXbjOmlgiVR34ENOmRUI6GbUI6OXJnTmCP6RvWJ
37aVEITTacd9IyBxcjx543V3jGSRMe4fTklfnYo46vAjV7b07cyOkCHVnoWo6TPF+8B/D4cJe/wb
1LYKUh0eWYya9NoBawc4h3BQ1wlBp7FLVmWdpDvHFnMwSxZ63R7vrsUb110tPqznFI9+rtzf/ac4
4/XRAdUnIwRCjRNVkEKKLdS+a66HgJVZv4CZ4agAGZqP+921YZTTw5WN3OtbjyKjTBFdM3NwzHXC
SN6c6EeBGtRTJaVdFD931N2fxJRuRxqVR7SV/FDNh/C2PbBemyO50mUHorWkhjsKqMbZxzAHrUtF
ZEHc5eBaeEEjzX5219X3cmlVSC7BG6w+WYsaiRc7/X6RBQwrjF/y24d5ymACon7qQwMdQXaH20yA
KaIKRzSR2c3p3dpn+0GSiabaLtkRxINMamr/OCvhN1xwiZ0spb9s2TseUp4eNHZPaRn9MMg3ERgy
rF3+CWA5WnNf9D0xBQDjTT2uACdVREuomXpqFkPnznDS+I4T/j2Z9tY7BIsuTfiq25ymMAcE89Fr
7Qu6YsOiehTaas7mtsbMcqY489xECFMWW2w8eY6tP6o29M0KHTHW005yLsdxiC5orwX656i3nZ7g
vvebizT+Z8ofr4j5sl/lWkwBGDG829YwUeaBo/6DwVjF5lt1id4gZeksAxlsDKHGz9eKnLJyR8vN
0XJ05uPoKp3zKXzJyMlB33VJbnGeTvR1Qo3Xlt460lNkAQj7tqatpv7E25xR5R3dLGlNBblVqbKS
e3mMO5I1Z+ON/FuBTsjWEBZTAMpuyeUW9c/kbbibeoK7SGOQIR/zYRmgVw6pMcZ2zQPXB7NmY0hQ
79v+2JO5TIR9g754V+ctn7uRbcLA2lYL+i/DJ9JOmvIQw7u4KxYKClXW4IhOkWBNhMHg/UAkhmBU
Jw5KYRPdGYqZA9w4o01DRrvSdgxcrHOgaslFIzmfTt2Yk6nUegIzOCXI2ni8+YXjO5UyVytrVKHS
J9A56GkzJIV6+q8L07IYFe2ehF1uKV22KDQ1mWWZQtlErTyq6yIRXMyvWl7Z2qB957Hny6/nYUbt
oTdoLfhl/jr5Oe1p9jhp+IE57O/kdeI6zksVzaZPmfUrL61J2cOKV1nefC+XhiF2FdbTHR2gFV5R
Esuy5EMG0y4KuL4jG8WUu72FkziaeW78QWNBo5Y25nSuqTJK/Z2HhR+f4N+Vz9QFBhG5h4EopyJ+
zp30T08oJqYyZo/Ivg+/kzDJy73i6s9ykQ+MjUXdk4p6K1RN8Uls1tChk9UmLvMSrKndQQzfz2Z4
9oqmlm/vYJuM5dXR5r0ksraAOB9nTY6UomcLR1fpCTdZdm1QeS4RxagSfafO8H+tqt8PvOYMwZ70
2A5muuiEyHWN5hnWhBp342jnZCHjTtNUhMCRK8duEV63QBRCkTFbhkSzeTRWSehecsxy1XD8u0am
TKH1v1e+WlzX1cypU3NPcBX0Pt8ib9rxyY1QSIX09XYAMHNM9H50c8PYw6VOdNahKTyJSDVvtfhp
UZ33d/Byy9s2g/zwqhb9muWmhqYLnGVE+pkSat0mA3iuxytnk2tpI2eoKEsk+bypvkexelbeONXp
+2r0/CH9w+0rb3PPrAm6uMf3OKUQJ5JDmL119JnBYyMChrRvKhr20czlSTkJadNifGSf21y/Hsuf
Cf3XoM7vN8K8E7q3gaOzCgnNSSvP7PbDlgh1J7mQusJ7rHYl0jNNWfBcfLv6Q/moN2/MLq3ashSe
is8cTEwT5OItyHGrioJADels0I+O68jUZxVrgulzi0Y0T6dlMHVAGoNmvCJ3gsxeWgNPqM2SNZvW
Xd8MXFaMbp/9r4s72qKrBNotUgvjYr0evL6YbBY21z5CtoXYpbCVRtzB8FtjlpdmqInJ9GI4BLXp
Ym2MJs5PI9LEbpbk9VYSkIrZRCdkA/sjqxgLmpataAARguq+XMj2bULygaa0ZJN6NJM6XQqf1rKH
NuunrEGGd0c1ZXUVSdV8u7G+dsjTYmh7CbzvI+SWiGrvkpEoBf14T8XWqSqn8D7AhIilWToDQKNK
vSMSUcKvCzcdlwlCEarHpWixiI44eV4IPOf3I68kCxOhw8E7B3HIDJcADuvU6dE8EdLkjP3gIgsa
C4ENd4xVrCpS0TEIvOqDvhJyVgRwF6rDsaSrYFgcK1pu77Y9Ua/tu9Yba3I6rozmQ1ty29R8wEzr
klsRw7L3z4u5sJrs5Xl1wVcDeHwvTDZ/pzhs8Lz/o+A7VQWt2A0Z+1Hk35o1O8o7JqS9nbAN5sRz
MCNDwbK00jznWVteuaWQC7nXjEz+T3uT854wqZHTCmqx1HcdLQ4myFmKbN/Xzc9WMa58n7+UqrYJ
4dN/oHfVa8hN2hLBIEzuP9KYHJ7afQt3MbW9U929FiO4fLEQ3vwO7kxeXNh0k2ek2c8hgXDnanya
L8CSNoKQEP9QP+qnveAd0+qioCt/5oXafUXmJpNXCKfgArNHJ5EQ3JcRjTsE/w1424O3PO61udlK
JqlI/dQ17bV4mH+PdWWxryUa8cW0lQEN895Te6ceRJRd/ZeLd5C07OWW0vRchNNTS+dXnS7c3ySk
R8oprZSNi38YKKKcM+5Y0AzWkC1zKL+WQWky/n6TfuO1bcefcU/GNPbzkb1IdTqFmOXV0XSM9Bnn
w6KvN5Bh24icZM35+xKJhbEe1TzzHQ2XxI30N+2zYfgwCMhRnb0GDRmm2NixoGyJEeBSQOm7xKf7
OugJ8FbaGmtP9jKX7bA+a7VLsS8bnsVaeKzOnH375+H07sARd1SmPVJ8aM8pzeQP7ap38ugrSbr+
qhUBqd98rzaWZel3Lrce4fAa/2xnOBA3hTpVgnHXxND3U9N41aFCD4sAEEi2FJSyDeu1Et+mBaZV
jNUKR0ctZebRfo7Ng2YRLCpgvnhPAJBuUVAPkCi/BHGFdWudgdxq3v1CVOxcth4sv/Iamb5awiSK
EzkpbcjAFPEG7LGKUh7YGkCpMHwd+xpnGgCIjAwbcgDLeQJxhWUSPEi6WEYZQDQ5Y8oeb/U54FxC
FfTe74ZPlOpdV8vSomEMfJwT/q0WgQluq2GmIdZ/OiRmyDNTALqQBl8Cdh7lOR2u+f7LT9hv4AYn
Yx1m+y4tUqfy4VmM+cG1ZzocfKz4nfo1tGDi6eID9FXnc2BxREmfZjJFaVvXxrQudwHIThVKXp9p
o9ZSJKPB+EIsbSHTL1i817N0tJmZdfel+sAxXlduDaGqVJ/gNwM+RAQUyrHmw1QH2UA0E5M55bdH
8oQyZ9wFevQjEdD1ECqhg8AkR4/5uqzJ1ADj5ltIv7hwd8VeeXM0YL+1kjOz26IOw0RzvoQ3kcx6
y7/BkGb/h37vwdvJmtLinWPb/h7O1LpmM4cUvSfkRLVhcvF1YKVQZ8DCwHYycmLxQ0GZW3IpbMB5
aGhe03UI8eh0ovDCJcM89tK73CczUbTtqzlVwcyQ0WRArDPkTaE8U0Kt/6QmJAqZNdcTip+ujBjr
JGxJ+NsvT9SAbWGTQGt6sTnEJ/X0tqhBXkMA8tqpFsJ6CJ1KN/V7YDNSQQg+SO8XYUyErc+M6S1v
3fBbuEDE8V4qhlzjPtEU/ZzQYednf7kLl1LAT8Cnaf1F9WXM3S6nbEQJC60F9FNUGynflp/txCb/
Vpv3dZxpUwFQXcFa8rRvtL+IwYhYOF/c155QiqPCdV1lHvDO+5uxZKM8uG1995T4I2ZKKSDGAN72
OSnaXhzv3SfiEwbMAbi1OSQh5xn8siMCiV1JIu94Ih/iiYAyoNXNbDe83H+L7DNA2+M/iUnmc2fq
VZnDsysYQ3904KX468CfwboOVjKKpqXM/emyIyECsZX/by3HdKjntoD/yG3dpVGuIvFKv8Ozepl5
zh+uWHMPTKUqlp7TukRhm7ZGCBPy2nfwREIIKI6VvT64bw3CFcIyQnYpmXy/c79XywZ8c43jGhG6
wqfE+XuR4SlR1riL1I3JUU5GhHgpYPxv8Lmgi5aKpq/8fE4dofFA40UzzJ7loAQF1+4REu41LhuW
kKgNxryoHl2AxDiqN9xxyVbaITlGBGqBPWV4Z+9J+g+R1gqEsv9ranoSgLmS8LJgULkQ6kPniMeH
tZHAsineREOUcOxx7TpbENTBvEJwKPP37pPEA7U7wWuyxqSkK4GA8OK6Kl6lBLg0mPfRoqiTC7++
mMSlpzR6negaQE9VVn28glPFFLDBgUIXjyrQNDwdgJqz/rfsA1OKD2Z8imNUsfOUi+hP4zRRVD2p
i+sZWZcsHqzIjKxxD3dZERUIdLbxmErS/kFILmOoykCtMelPedW710tP00SfkrzqQJm0QRZh9hy6
0t6ku8jUbSr0gWY6M5eghoI0X997pFroHq2pNjEipbIyvK8tt60ENAD9QdFnZ3RUayXgdlOrB8NL
p0LFjeZl6AqriQ3+9nqdqowu8frm6prEKtVdlAfchEvUksGU4jr+bDN8VebwOtPO04mKNzHtI8QA
GorkTjuDBwwAH6ZHoEEX42wG0c1hGs55zPo1+DQncrT8Hpnnyu1JiFDu4K64tXde1/OMC5czZKIT
T+dQhm/LzFRTyHVx4GqE6IG6+Z3AmNeRoY7vadKiTHmV7PZLgibQlt+s16mE7uBFDpw0chMygizx
n2VInxnlUELKqIRENJVKHdaieO0lS+nS5x56x8P0ChDfJqInTyYoNbiUyEri23s6dohWMvL47RXr
8YxZbxpi3RgUV9OesBFK3y1ucIb6G6s3Zf/l+nx9aA1NbRrovsKZGd8n/NNVKIUILzFCGIYTn7CG
+NWWPGPXAEq0nwWIgFL+hbC9xRNqLdxjxOMho85d0S5q2A5q4+knOqIg/U4/VqmLlXpius56HVaE
LvYwRsZGssEDiNzHiEBch5puPR8dGAXNYRoQIsi0JaddL5MbaCzC+5uQzhD8Xd0ySVo9gZjNE+2Q
cIUr74iN2fomw4KkgDoQIxSOis4r1LLs0OK7zz7J4SoxV4VJx/fzNqiZPk3ZnpjM2l2tcvv1DXqI
9vqeh+DSa+88dl2jcIGxAKrlhrttzf0ltBs6MM3oRt9cUm+G7H8wVlCc6S0fVgc2R7WuNX4O3YVp
APap4NL0l0zWvelpLcaKRztG4lwZlvA3vTIB+utAV1Gs5D4Bzy86HLgnLyjMHsCqxwDj8UWhbLD3
fc1hLiKQPyjA5jVrc0Lu2zwjHcktbMWbsB7WPXibPm/yfVP61DR322DkKFeFtczhJJdWK4i+TmKd
e+lGLrCdKnWks5+FrltL1mfvw+ytaav3baGso9ZBT5EkpB9l7DWNoAazxlbbLRouFui8+GfJguu2
sIIdZguhduq7M5UecfY94Q/HT21d2zDpq0EXnDMZxdmB96iu39nhyPIz9XMPYCbixXudc2YgZ1KT
9/1MBpTXd/15PGmRDoaAR9XaVIi69A8HKWHBirlHBQ1ORj4qVZ801gjZvwyl59OX2LtAcwDfTvcb
wGI4WDlUtIsq8RSR2DrHG3sq4mYGircSHO4KeRf4zhMvMifVHu8KayIuDa8ADeIPOu3FM7GepHJ7
kbmrA5YDnfLmmxM2CqE0gyPlRwvByrcFwvDWkmVipJZQO+zsyI/62Ug4lcvZL6AnEwHoxiO0A4rY
djKzDSutVFx8xI5x5+1smkbpRHV7Fqw1EnudrNLB4WRTJ6sc3191XxqAyA/TaLU7Uh7+MWB4+u62
0P83jCkKg1dhb22vUn/HGqCPBMCdkIXzI8AEJtLyly6DpSwmRgMyzVLS29GUFsKgy4LYztibF2hO
utqFV3gkgjIg6Lj+2QRExyeWskbpzmqEwtWdtAJLHPyiwvG56AdLiwKG/C8aFNqfszVsOYBsfqxC
B8LI6paMvqGpBrJvoyAM8bPyoCQ8TcQFai/VYCmJAfcOmCPFU1M4zFwXIxywU3O9SifDMXIGU9e9
FGonzGxWCuDaSB0h9CzDdwDzzM/XXVW3b4hwLB/9Kr4KNAwlpI7gK94jgoGAgeJ5pDennwcscqn5
/9o79p7/lvlDrgfkAtaQZETsCijC8t0zO2KVLur3kDxoWyoz3LnQ2N2Fayih6/vJHp6JjwLHXMmQ
K6W6pTwDfnIdtbNnInx05lUHY+VwGQ6w+EJxAyGufTPbWvtBilwUDVBcK73j0N2fkz1w8D49JJ6F
7vSbHFlp2IOvnuD4oRwzstoNTNZQUSeAwZXGi4CKj32IxZEs52bvxGZOkivkDay9eHDaHoKZ6pOI
AC1Nf/3bRX0J0y6+JsspCn3Dtr5axLRGtScAYjMBl19BglSgV/Bth0KGydsOqBw6YRtWJGXh6nsB
6TQ+6kcNdctP1DfT3ALStk+ZjteAuMak/FWT1aSGUSvz3EVjnKjDbubZVmX6hkyukBXZsmUDZy6t
tDpXc++o+Nhgdy8wtgggkhz12DSYQhLNrQ7elLR6zKea5nyGSLJFKT89CqD7QnrbCOoNLtTfkk71
JszUxZJQgTJG6MukKbZekf2fSsfxYxPHVVADVpeTordecqd+UCQm8qMwWo/KJHuqDTi6omIMpENT
Azvb0Y2j0LTjDClA+amsDgMnBnpW+dGxNc9eAwl91GZHey5QaYLWCNBKKFw2LghldgMvbQSSsjfk
tqmaxvEnycVMEtLxnUx3wtUy1XqghMFgXgCxJ+JsM+PHvKoTVav+Ya0zoZNUSgZDfP+Kh49qYYyk
hM6s4hGQ39t8LY9FVQi6VoUB10xEYS6fpSdn6XgsLLEIZv7PSrLBth190in7Ce/Dd9Pp8wWt/Grd
iqcEI/4+bvr6Y6/AaM/KFpCq6i0t+jG43cqzF5s3yH26bX8hqJi4Yklgfw6YRPYbDIYpJp2GkbnK
tmWnP0huw1oJ/fN0TQMcyDkYWFglKSH66louaHqCS6ogjMjJ+HgfWaZaCyM3NjHiezNzPUK4NvXe
F8u/0MbbPGObtKucRlQPoDuzkrxBXaI3SjDqNJZtMHAQ43hsLaIf86llRZiKCLunMX9kcrXSsoVG
SRF59S48HWwg00vSFGRUylwqnOb4u+yNxYby9CfCS9P3R9+MfdY9sLZKmTj2tYxtT+rS7znD+QKy
AoiHZgPzi+wlkVh98oPwQ7QdjAI9fxQNSZ8AtEYYnei9y3uTcPZ8VuK2uxOorIGRj5Jb8+6QtffW
Oq8EVpwVkK36+NYl2IfsAJxW6oTj2hysygwRXLQB01gJOmpnypInQ9YK+2A/AgO3J99tA9vaubAP
yv6fnCy64ZIldQQZ7TDbukqX8T8pn3xuP2oo1nLFJeP/TjWMNKTLtO0AMmPAJka/VrIAmkX3rWVt
vcjDlzt0FJVOWnxHnpm6rZQJofxKpby/83C7oDYx2yMIoDapBhOQ61tb0mIhAzqbWWbOOt4t3SgP
qjqc04QrbliBPXQ6ic2PVhy3zfcqgX7zxRJ3V0dMvxi3IRziBJCvpCGX90wBsGey2sIb9rmBLPV1
rf6HLOtBrXb6u5tMLADC40TQvFYvV9v5CDURcc+MFoliYcMQL7dg7Q0PKI304mf24WV+keTuvqCp
fVqWL5kQfzRTLBcfHit4zNt/EuBLQ2JDAf+8C8s9qYXezHrvlzLIwcWbCuXoxdGjnmgnCccSRcRP
BujkX0zHvOkC9OcqhIisYtoR/OF/eJLZC4VSZUfonen/t2vyeMTPskQ3w+C01zfssxxJJNkMRkXw
wVqwpIyQSSfeBfE0i5Nw4gedb/GHoUVKu9m07Zlaqurr3OZPC1ggjDWXfB2E7Xs4qKmkKCsQTk2W
9g1BHqFbicIe3C89Z8vha1Pgq44yyUzaIobdFaIsivHJCRFy29+ZmwDd1Ytv+a31dlpFGQAHz1Fo
shRYLdbJ4EPxVUxzbVSo/FElSFWAQpp+y04Em3sD34+XrI4uzBWUXn9Ao2ALdpKl6KF/k6EMXEZJ
8RpzYtQLepKUOsvA/SEXhxpNiIiVuQsvOo3RXz5rhUB4oDW98e42MWsg7MquyTXIico1RI/TLsBl
qkPwPKKPXcv6FeIL7pbBAQaHrOFuwOv9t2gpXwo3FI6JxwLpEYMvhNaOxTy0b5xjiV69NcvzaAcu
aUzYYTgzo2fLLhqJahrB9cSFzZ/Bo9Z1gPNKiGC4dWF2bRmnqDiL6QB3yjj9iLQEqWc6nm7hn4vT
sMEiBF8LygPf4P6JyLV6WyVUXxjcC9qHLCOqQszFhNUebB6JOR0GV1SJo7jpYHhBDsARl+VsVYEf
L6UU03o2V3kZkl9ElaYb9wULBwkZD/o9pDsTrsuYKzBtTmeJ9ZwhqW+wZ/M0nd/mg4q3UnFH5Brj
5/nfZnve1fOJCY2OQr1rFCW65W3XFFgqfGwkF+bX5TEpewFxh39/IthTbp5RMcHhhu+rLNQbuGG/
oRDw+bybBtowY0Jus45JRRN8/zLWVcrJdMTuNb6gz1e+oRfjICGZrGxURPweYweccQe4C11tBzRu
br6SNO4aUa7gMlxnDZoQ7I4Tq34ZfsP7HxiqG3yyGsq9uarfUIB3BjuLnIEK5RdeBoJ0+kVDPI4K
M7xBsdL3nVyuA7LrASNM5VaBoplRMB4k/WvGydIkMsnTk1YdU6i7w+N9Bmj0gTDdK6jyxILPgpg9
Lub6WERXXNgCYwGObnyPM/Hu8YhRaG2RrUMX7Cipxlhx3oeK7/7n02nJfA9Uvc/tv+ss1WsJY4ud
I8c8yE0f6U6+dZHrECrbuLM8wQh+CtP6rDOs+dwFSdhEVxAVHZiMaDLLP5MGfecFHmCbZF44K/+B
UNuGcSZldqe4WYEEHFW/qvBkjBbREoAWiUEgrdJ2rylBZOY8lAeYusaKM1UErFr186HwN3N/1m8y
NlSrWzaGTdL0DyhzvUBGpT1UHCTsBtbHyrgl94HqfD8TweZR9kFUtFuEoLsfl0VRSXlzm1nsijNv
yjtdF7ZqzPUyxKZUGkfA0oDtHFkeFHdvR2W48yI98iH+8/XC/R5I1yTrq5y/AH4FZSVwaznc03nR
AebrSMeke2bQkOXuPwy7qLW+ZJSuouV8iz6SlN+/2ss0IHHPgPTjHhKsxV+2i9Oi4YvIgBNYcdOD
CB6U2vqTc58oKKi8xo0F5cXU5vGt3uiM3aju3TUYQgBJoJJP7NZiveivBzEdhlCjJne5ECDHMPly
xCtY3/sQW6dF+Jy/QGdySL4jxGcWwJS6WggsjyyNIysqTsw0MUbDhxSYx8HG5k3RJH1Bs843Z5YW
EGMRz0SKU/jul4vKymDugQiiqCBKz6RQryusir9usaHga769E/SsqCsVcm4f3Oqg+EYqAFRCFPbV
1Yrc+2TmexN9DFgtDvGxyVUP6MSmx1bs1TiPWEicEB1Fh1zBEX3kT6I8POnY6x6cGuaLqbjf7nbR
j5ydzw9AiWHEoPfvIBzCZYSupyqNdPkZCw5U5z9SNUaC46+Amfg0al6pLjRu/nAnzDcBuMF0vk6E
0PmLQqc7WtD7kaTYafIYjIUkDVApWWFcPY4UI4mWeRLBgZUR/AZgd4USzv/paZw16jv2au3qoAds
a0eCIkPc+D2T2TWMBlQPbgBeQphHt7vZQokhTT3ahhr6P8vQi3d32jk4XiUoiPD/oQqhjXm5CKeU
GIyTPU+v/N/zhwpl89m+1kEMH1M82fbz+XPy0V7uMe9Bt7rxeJKFVSWRGh7v+XBLrY6DHR7YMFfO
/V1/7z25S6IIhPAygxvp+AflvNw4mtMzXJJs6zvMTeKkQ+hf+Pywj/DU8WU4JCPkY7PpCJX/TnRA
9+ZB+t33BtLSLuIZk+V1qpcY6JuBfn3HuJHuHwE4BphFKUuyp/77jTKXnvl+El4Cr47Au1ifPgyt
ZFrWUgsNunUstkXDu6OtFUUoSblam1rPipsUUuakUqa3GX10XIQEpuxTS7Kfzw3EW1Spl8kvQXkD
643g5zuwQ3gB+1eSbI3J40Qhcx/4K4Rl7tuUn/yrTUFUD3hCjNWu7jrpQzgqhXJjSKfilMuMfElv
qbn2atRPFR0YaLFCcCWGtXSX2MAygquay1ZximMkfoERyZo2e4PU33X2GUEAoXyzXGxTEAfN1u1K
NwXkwamdbZDNXxI7blQ7o7M+TBVCJSgjIAMJRIHJkSBDnnNLZzuPXoREBdIwjmRodsg8oz4R+kKo
xC2T/srdp1vGP0+N93CSBvWeLLbXrcQZ2aIAqXRv81TuYm2rMeNhNw6k0u2P/Knzc/gdQvGhV/sS
7GCrDas3SbaJ+qSHfrNRq6/IwDXDWKUMDb8bHWWgXpePGV2XPgvHrEV4Ln3XEWmI4NTs1RhfX63E
U/21XuMCa25ZzXpDhP4V6kZnd51j5oCRUgPYz9fn8dhI07jjfatUC8cZV7thBhGVMOWWzCo8NELx
ESnTlxnF1QF8dWsIe338oVCHXJjalF/95u86mOXLoU474NqUdzjfrhVQhCraH4eHuDI+A2HybI6o
vg1KF1wFmQ27aP3DPXRUirmprmV48hqWuumVQrYS5WnCeKafdsOnn8+PDxnfuR2kwsAcfzZCDUPM
jbLI72FUqc8swAPKt9R7y3Ch0IYoeorXH5oTnFIYhj2IoUpIbqGSPzyJqBzSvwJ/kNfxzpmykfGD
Pt0SPJHBuvDrheBqgROMhZnEdGbWQC1Ao0K8wMJEhMj481TE4BdCPhntFNq4jZDLFN+vrc5PorV5
y2h9/rgvyUomPFcfAUuXw46QtFiO1loGULDcOAL0vRU1q8lrGdy/P7Oml8RmrY6SyCdIj6W3Yr4n
PtWB0bZ4PFHNNRVcfUbPueW4RlH93z0edIrbFL7Ao07hdPKKpT4TZuhQFtmU5fc8COGG9grVMql+
pF6Kl1a9CwyoaCfnrFKAAm+tCETOTJ9Pmm4+Xld7tjtL1AuFyVlwgTIt+XLjdv8dtF8axAkb9tyK
D16RVHmWzBSuDmdEN6xxJvIzvLpTfw0D9y3NrHHRKEsLj2HSDhaUuYGDipaKacc4WWUypKvcStE2
Gn3gzoIkvBSoAnBN86TtTMBjx2JzxWZddP59kvca7CpGqDFBKOMSXTJgQf20zMlMUBwVGZOPdQEB
C7O1rlhSAoEQlORUrbxmkA+uJIOrxBJn+1z46XQ6ndmq6Vjuz5wKsO/wDCxIQU3OZb46aRsHdqzd
2lMabsCUFlAFttlWaNcTZ3AYeFSLH19vozNTqEaNsOY4J0/a97BPypPzqGG2xr1oyO7rhBIxADOM
2fHRRa89Kf7mgdqs8Xvc9xdyWOsgeMEtqva5r6WBM8IM/2WiB4JEkt3anW61g2uMyigpdiM6s/4T
tZZLPIXEhY/iwKCbKTyyPkJ9GjzcYfdYppBRr1uaAQqj2/CN5AP1sihgQYEi+qC77gzdTQLnQdBz
hIbjdETaOXSuto6oBwFvy4QpLBwq8Rgzrgfe0qJkHTBryPNuCp8ZqOYI0hkB3c4LE5GV7R1W5luW
qTVHgxvcr65zkzVY1JLAUmaZL+GLOMkG/CrbkTpXNlsUK3PvS6eyHdx07VDMKqt4czytRH55kQ7t
BkNGL04uqSkE9iGoozJfTZQjafQ7LaDPm/NBXuWP39QhqSfRAiIVWqcTwf94RhPNw+yxQy8NRO2r
M5k+qxa/3sgBqMOpAp4D4f9pmqLemwvv0iXqu+om4q3sdGcq1J7tVLgGyDOJNMFhz+NZ3mvj99zV
t3QnhEEECTUncl1YKIWCZDyunNIvl6XNc+YJyQayiVljQsW6VUibuIV8dkpWLqoQx5wZ1X0AM3SM
PEshOgHIsFVP3ozrB96s0e8k4Zcu8JEIS7Prr2nHzB4uYQERwUxfZeMDBN+ZwQbfxYsidf7u8P3W
x0PvVb33I6WDppFDo4IPXyhbCaJFfZ86847U//ZRopYd03L1yLmkf26xvk5lmph+QFYXWKj1cKCf
5zj+BrgopBkkz0z/w72u70+OASzMqpZblMY0KyHumuerCaz3RFPYvir+4Vu/9N9IKCdiGJhIzcmZ
7ndt9BQH+GI4hhuEt+QQBRGy+mPtyy/20SYoaccakVo2k5DPCKyKUQlT783NMpxaJBD3r8vp0Yaq
XJTCWBvK36LipfvH+xRa3gPUVSK5VrFbKhm/TCOnNu7EGkCdafOC4Am00Q0egt4WY9TpQ44piPg1
wsrumxtUodtTbvr7jYOfz8o4RaNVwOE/ns0XbjDFHb0+GmOGHhsqTxZy8tAnbxBeUeAZ36oDo1zz
5z7mhcGeVwHIMlWDQIzda/iCjKLs2dXfkYh1Xiq2fiBO4K7s9yKDkYwDsnRLkSl705f70A/cJm6R
gfXRZMSG+amI/Yu839TR4fo+KYX253mFpotA7/3M9CdKvnV8Q8WeIWUI9f8DwnZ0bCQTzFMMD3cs
uOLdUgM38fOPum4M2j+QYF6Oyi6kcWQun7JwxBmR+wMm+DmDz6m1O+IoC6MzKXeXtd/9tay8QaNF
z5CilSi+jI0gLsdY6OXdcwhX3VX+ntrBNvzvEP5nBCAx8MdGrq1HWHI+Ttj52V7xGEAyNc68/iai
cPsRFK+oyHHuvoK2z/h7jQw0/7y10J5R8KTFikexkvmUVhzcoyjRGVa3uzX6QWxlpkTBQ7J4NqHI
pyFj9z2qkakcj6QQa2SCBgvMdHG1sSo+UenMwcUcJuDzj9IFbx1ohb4vCVM0q7IcSTb+Mp0Sy6s9
5St2sxMittQ2SBY19D9cFT9HQwrrytJIJHpIvKL3xkqaQVcC7zK7xRafyxOaTdo9KALgnj5Sx2Sm
lF5wIeCcX7aRlXwStlrpFLRKwU7Me4kksdsLYnlDGd5Wsu25CRBVxWzHCvTNIUBa2bIw//kxJZS2
Xe0xR5cJ2/VE1q4X33cajtg2bh304iKi2tSr3PfTtHl52NM4ICgnX6IhRhePBmdMlFv2XrHdAOwj
SIEPEs8Lbon5NUIGt0duDN4Iq9Nc0nDKrOjASlaEvNsRHd86P0lv+6mlwFuFfTTKRxb0MWlvqmCb
3FBavxc6tYixkqEv1aiioCkNIrr09FxNKDDcfAYG7Zja5/gjLK2TAxMLjpYrowtYfOi0c8C/NXmz
4KhVIOb7JpzlK7UQQD1HWIcgBu52VrSbDsh5N9BO95ZM9uM00Jd6yeM4ezsRlgqjyb0uh9uuhjii
PvNum18N9m8s0qjUqGeXxw3IavIEKr2lqbYz0wmpAmzkFegHP2ZBonpY4D6FRip87gwJlozvA6hf
9TupVKmdl2KctGuZL7RhGZVmHJuPGT5FzOPO4lic7Idy6nq98y0dPyVNCSYa5d9FoE5NloNAFlbn
Up+2WhKLuKP0kP2z1j1ae3eK9ZSx381YnL+Hxb5U/JeU4V+/IWdTx/1uTjJNG6ifEw1BhzR9I3pJ
t83RZ/Kbg2ALdE3t/A+QUrFZRV/tZbzXrJvU1S7trcR+OJ7NUP+dzuj4dmTQ5yf0qbAkSR/c6Pf9
CKuAxUx458J0NKvIJ3np0uReXvV1KrmMxJjUJDiYIeqT6za+WBf8bOoRjKEXdvHiu0Eir46gAK55
WXnlh4yB3i0r0//sA1hJYiTsrXJ/u6Tinu1L0anDdGepmhdGzD8+kzG6zUzc3ZczPgALksjz92Ha
NoZhGa0XQhJZsPYtfw8U2WdEHJoeGr0TGYX7PXl5VgIfgReKLv6HPEg6Vl2e3PG/pV2zz+XYbxyw
ZTzuO+EDxY8LuxvjFJ0zvjDr4dU+S2WmfHJqNqsixZYdJt73Vj2iRRZ0hytf6HyF8ydWqQY2M38a
M+Elo9Ob+gxKS9YOJpFiuH2xYA+rvjTltIwn7CQmhYXmg5BQ5h13+epAF191GmMHX8hInP7Iyev5
GScBmZOv16cMVmdYb4kVY9ZhyxCQ/3IlUkS6vvDaQXH16K5K2vLpUJPDtI6rr/NcGZXQJp121vk7
pBNcTg+wrwu4dQsqcgDWNqkV5F+jiKC9NpYq49Rn1qQhSrKjFpq15U8cLsTl6MMwWKLuudyPZcxT
vnH6ZOeknRvegPe//wIso0OLU5Roo4u5CN/YWH/krDEd8BdV1WPeDRAlQnvMgVrNEjxXKgvi3YCt
E+GOKOhnUTagl5lopLdb+moWvJ3uv0/cR/ZjRUfdyMutvku2f2Sz7B1/Cj8zRhMxeYH8qUma5nEV
AvkCVreH6Z2bFPpa7HopkBvU8ktIjNfUHYEYmmk8WdiJw0ZyGmvlSUpQC3cMCOQhkedif5ooJiVg
RLE59znotY6+Em2/VIfDN/iVOYcbO7iZFIRToGmTB4PeutLEmcpWhSb/TQDjx+r6/NZ8KdODDQFb
yGA7+LrTtVTvboIkmgX84jdnG3Rj0nuFarFQ8g30OtT4Qc5sceW0iyqJadYKzVMNLgIiT2ktYsgj
LhJOswBV/cbhXG0pvEH169vNWg2bLjyOw3nVU80AYt7S5RD1VLxHwO2OtGJC4AEuh1h2/2Owwrlj
C/trlbdpwJWZplUQSXQnQLC6OzxgscGUbvlOlDI3WnAobk3yQ4XD6snCERAb+WA2hETmVXWhVQXy
+4jsjHFs3zzlJvanyAkjHFQR1SiiGfWP+0Fhnxsf998aeTzPvomXD/k7pYmKL/T+1Yy0wP+uKKkO
qjrG6C/2cm/GN8ehcsfGbc82E6ROinbOoDfK4RS/nSzFH9MGO1n836/YIinWe22JkcT8ilkEzSe2
G4fNSh7vg6rrygIHcZg6vEU1bH1hixu+aOTVkbI7+OP9doz1mi9UIv2sPKMdthtDodBweafmWgur
Q9231aS03Gcn7GqSXzYBz4FAYjVzXWvBpPj58FxwPuSs2kN7gORkWtLrGYSDB9hv7N33xZtgd2JS
ejq4q169YKhsJSEXM//PLbOUGdDdQtxc3JrR6X+hthoWN6/ND6SYjOvPVAJOHqLF31LNumD07XVw
MmmQCuUZd7r4LQIG6AOxoOuj09zzwvAfiOCMkiqDNFy3nGCD6kzQLP1iok7MBLhMyaSCIQ3WmgPX
uKMBuBDNLpUwyzAxAcyQYXuvt+GIk96xRf6JoGZqVwamrSSnYdaK+cugcKwO2IadEwObjOozc2Cs
qaPd7+XHHEaWO1tappIz/a/jxHHjs02E6jfhbJ+yKYJPXPiqNnvpcAce3GguQT3thmL7yNiMIEuu
y5Tg/kdE3H4r1hHW0HliRkzwvXH9bQWHk2JuLKCtpgYDQp2wENRw//aLlpiCAFvgv4P8sEq9qooi
q5UmgzJx6sLCeH+pl5hpw0P+ZBx1l58s0imxKXl6+kEcKk+AMhV7gElfbMEP/yYfk6SDJHWIQ8am
Ae97FERKVaq0TOOQUXVW2eHAFLwZcKxaFYnFhDed2t61rgFM4uaUYJcmOEf13d3UM88cMWKYqsyz
RbGhHvxJ8oSNxwjwbwH9Hs1EuP48G/yqiWDy8de9BWXxMNAEnMed6IRmUx7J2fAfmlHC0n5eSpVM
PHGDaSxe9pxafjkCRYGNZq3hvMif/SIN2+e5us6So1v+q9QecfN0Ba8tgoUyhnrxVrxZrXfQF7HE
4c+G30IN2JCxE5duOCe+oKbcig1EddZB0h6PBNTwX542L+LnomeGMZd4xekRHy8hloeFkw/BDpmo
NGaC9M6g9+U/FcTxVwqhJY9sN+wsn0BrB79L/AGqjfBi8XexFiICWi2Zi/3HhhxObT7VsZdhgAxM
yYzOFLaC8kufBHGfejOs6fAX52fUXvZvHs7sisrrSfMjf1yphu+XJHALhrsCQR66WRJ3+1H2WY6I
/yflRm0MRlIcPDbFb5ogf8LXJD5Wp875hg64Da4LZtJ9JG9taLfAe9PjMEsuxxSpj4GJe8QB6qoj
wvB57OZq0SLfv3RhFG6pPSdfe0lBK5Vq8bZdc4egexcQ9D/dCLRqP1Xetv9bt8ww+qPRBRfAUwds
GlbyoNQkwR3NYAwx8QIV8XCKX3NRaLvDA85+Pnv9heXbxgLpaCb8B9ntPO1Q5ch4atZ59/ZFJDWT
nmwjXgHbc+3wVPkWImA2Af3wn4xy63/Cldy9bjrPll4C0u+QStUsvy0UNxsKLZuhcW7UeC0e/seE
6vnD0M4d9z9FOSDBP46n8NuUQdYcRCoSjT7hrcsalMdtJrl3+YuH416s8Id3Nb3CrQcN/56FEw1c
AEMskIbivgv3R51BBEGVlsgTxya78PHxUk7wG39I/u1Tpj4hVN9M273FeE6ZghGLdDvrAmiXmY0e
tmAyulEICjNp+sNGH4D/naFSqcNlysAyVXH7uQw+m/h+aYcyDXOHIsa3aqrW4iyjVOmZd4hMXbV8
BM1sG4qbGwOZXOlBGHhuy9UZhObf6BA7jA/VcbF/NN/B+9f3B6BJchEk+9Im4/qvNbhK0OCkye4D
XF4yqAepPxgdxxLHZ0UkTLppmsurXuNNj2m4sSY5tiOsgQcCZ1xaa2SQdbVqoJ93xWJ1Vy5Wl8CP
LPg0hRhuKOeOfOQtJi48hf55NuL1+FkFHvAylXXl4DTHwPCcHIDzisk+Mo2LSAVMYgi7FN8ZODEX
sMBSDPEpGLR+M95EoE4+pnaDW46wowITrWWfWi5NSIrs4aVzzX3Re5J6lXIvAEIpGBMPXz8h/mUj
2NEUcb4rnhXujkWOLPZ1tGp9qjK47L59DJ+ldP0ThSiG5yos4anHSSYrgW1KJqXLEdO9s203mCIZ
Jj6RAENmRLKgcSSeojCoPZlOE9upQYkn7t5ZDq3QkgfZLntXKWCjwDCGcWubpnIF88v3aJyNkO5O
I05RZQ9uRApDoK8OcIlX4jmUTTrmrIbwr8nSNZ80BKn82IAs83ywfoKu9b6jbuyQxpw2PHeVA0tm
AyDf8x7nbUYLnPqGcEAFOpuSQnfWbweeyJcQ4Er+ey6hVHo9gQCMdDg5n/L7tGKM+Wj7cD1Mt4kf
905jqrgX4Taispuinm4UId6AWQf9NtdDuNnbImyvfOK9uHELxQFDlI0SLMTmvrYX77y7MNY5slkD
DezMzSvrc4gZjEJP2Sg4MMMf/KKjBnlFSt9MWxwQeC9g/8calGUkaExIfS70pGTXl0IanfUxy/Qr
osQBYhlSRleftCMpRbVANqnRC20Z5QSH7cp7uj9n1aTbxMkvl0AkjarzMHuDyvkzRpRgYWRZzVdH
Dv7W9vQ+He29+P6//Y4jgyoIb+ue9YJ8BiQfT9SmMQ7tdakMETRS72CQ5llEywgvFixXqhagWSZA
UzvCDq0Ld9pYCq5cZ/qYjFfGtHyq0PsxGYLT38jNmekk6cnSzh4pgCKBXzlVJtjhNl2w47W0zKmt
8HOlbtkU+FjBFKV4srw+6bw06lKUzXvx1z7oAOCm9u17b0mvkfZKtOa9EfsZ7syEz0MiEjd3ik4B
WP+pnOTCJVbIXq2FAzYj7zW4cpo5TGpnLROgR8b3JdrbONhFDvU4CRY8oE8Gfijr/nC09Q3Qp4FN
mUH5yjWLQBEWDZVpmSMoi4V02X8jtl7iLsd3tSjvfAxjvB68s8rrRUgxDh+aqdlHPhTPmEe3zKsK
wLzV66VRURPdJiCD1cIm30U/zDZrPxzyuOExIRX26B0wKHKqifdR54RXjL9cvHEX4NADp/GRr/Nc
o+6Lrpq/XL44CVheWazOz7m6WyT9YQxlt8yTqnyn9cTBCrALikX+yH4Lenenhy4zPKwalweSFzcj
7fFR4hNlpNWK07kWggjjFrfdvotSbNrY2JQRQuUmPcoEMLQL7HgrwFA1ZW2OE2M1N7Eq7SbDIF4g
Gqz/FMbXmy4TUlM6//DFwlxTGyxO9J2r4ssnWbWeCoYoknWX5TlKvlm4SEqtTJV8Gu4G/3fDipew
MQwCOHS2bg8FYa/QaSrDRU/9vdRw5nax1DoYQhM/tdIvO9ht7lupuO7aBts82AgEGXknJh0o1TS7
C+5A10uluPmXz3D0iFhmQ+MngkYMbJnpvu4Tk8964qxA6GPgccmw9q9ZubYnieF0uNbO8TFixuAJ
lk3EYcYr3dKo2nroTWYYWDT6OKGMGFGEkd87DKOe5pg41Nmm4Ictx/ugGBb+UWjD6VjRV2utrW+r
eqhXJVfEEpMM2KSS1brUgM24D+MRw7HtWa1f7S8LjLkN0UdNf9C58TzQ9GXvjIoR/4on9Oi33b6q
f2yFm1h81govKBCyPtgQhKkiYXYZaVF0wPCOJOcSK0PgyWgfBvdZYZCKE/wHuJKJwcIiDr8fEEaw
axiqYqVBjEe4yJmuZlM5eOKftmflfSNmkXr3x+9IrqAtYpfwaB9Yv0RFZYwODfN9nkSkKL0ZM2lJ
hIAyVPRiq16WMdsWdBJxQh4YLd8S6h1P0sfHH0iML1g0MWMlCcJRbpVupPYNihEtbJrXP9t+5h2q
2kHIGk49E/jBIcU8jwVo4bAqdwmCAiFlAq/MhWYTAJ8LFses0p5iQb25bzDWDlhAJHL2SSamzKJu
n1Auhd0YbyMfKIvYtQsdrgewBBfAZYI6wWBTvXrrIqmxcbb96JEQSciWjgCWqlN8Pr7YTmglCZLU
7cvVdyy4dRKgEYmHJNmqy5yhiD2/erbAtHv2MC/YXHquxsisdyylD44GpeqBim4TLk2YbR7B0xbn
uHCeY3oI6e1YbcOBkemfV6y59RwEYELlsUvVDCQkDtfsA6c9CfBgwMAmBZxFYTshKAkAakeSlegW
vSTH4r8XNicQMD55QpdaOy/skPxnTxS53+L/2UGXTDxUBBkGmpFmw79L3rAMhwIImPLIxSd4ulV7
016a3smRfudQrJvt3t1Db6XF52U3fUXSjaQtPRP/AbrB6FULEa1EwT9GaOqHhhdSPmKjl2Slhqtk
cGJYqX6Fh+cpIKGg44JzAZGEHk7+ayK4xUTzEEcD5cbFr4fUKLnPjcRVGveIas1CvcvkBevBFodu
6R2TY+jLpR3Ir94NfQrCeL2fRr6KqIy16mzBDGw73614DAcDjkX8CZEFpiYvqq59SKqH1ZKz5aO3
/mYxKK60U/ziFNSiZk6tbeOE8UcU3E40fThKr5XOrBJWrgpWmFCo1InlAV0YCid9LJ2pHDNOgFGa
TCWqI46eoBetdQFJvwTOU4eShLoaRZBOoX8QAaXciy0d8XxDN4UjOQGmdPSWllD8va7iepf/11Fg
c4Jvg4WKPuEJ9oOJ6qjMRLQIv1Gelk0eUfPMQ+HNVi0ihCN4zgyaPK6coxZF5difza+NRH0z+PBZ
kNYjqhuHRX2rjD9DZz67ClaE/7OHcwlGJJjUv+LT5TK2tT+FB3SomEu+OQvjiSBSLi9SEC5abiCg
ZnoIer0nx1vOj7O7rGDtre92yVRwyju7axCzWka12f2XrXTF7mRxcrlcTD9/lwi1aDP5wa6z/5Bo
BL9MV/a6TPM45QBWy46Wk9W9wCKmwdlhSIkaHeDSg4XvM/WmPF/1WwzIovOqKpEYTWzL2jrvI6eh
cjgQc9USMptS+LFoepDu+P9utwbk8f8NDgVqc71nGvLkoS4+n2jnhiaKDdmm19yZtvRKyIW4QOlg
Lfu4p4v3922/tcSBCoBcZEBifY0E4Vx4WW88gK7on//LNhwtAiA/s78t8vySw0fS4fDa17BDT1/e
gYN6zhMs3l034KW565zdwo/yzn3qWYZZEJFNBbc4k75btIAylpOzf0Fiixs2iklqvBnqk7P/vgcw
D2ScwzGiZp5G6n3XTgFI6l/zrFLdKxPYeBKf+FQURDNqvhpO0o2O/WKJdl8FWupxAfE2wNUrPihZ
wiyMDceUGSsnFlA2MMfC7q4QHH5rSKE0W9UU4Rk9TkS3Wzvof+cK/A7mvUrysokNBTYgqGdOib74
2z0SrxLg7fO7VCIAmOuIZXCyvF550bGDm0emkK15SYR4pqUFSSGfALidWEOvBtT/c5//w+IbJzA7
+AkmO5+hybg++iuY85Ewvwpk98oZ8O9JqmGj/iL0M0RGPyIfbzO8gbEUpJda3VsFsSmd049bcn+A
CKtrEpmJxmG3klGVT+5+Wm4M2fdCWtvmsTh3Bdjj2EN2esCUDHn7AGmHD55hkBwXe+KNoTr23Xns
83VIto1RdkxntHpg2FueXFD2rt4FRvxSvZgt5FTZSNgrTAE3XDjf/GNykECYdU0+aWAvou3/g3zv
vtmYh7t/sIhf3O1wNldtrmIe2jQCqQ+GD+MLypJRE61XK4oU2mhRF3TWXeeT5SdhOamLn2jxEhXN
WoQrNz8mFULxasl0uGuttZHiihj1XrZnrKWNjibA0pOvohU2tzPYrumvHfyuWbc8O9QESLgv270i
6w8SIwDc7/ZrLfLn/98Q6N4aNro5rFzlLqNqJ3EJFvJl3NYXu44ccF6OFtPiu7jlY6VmJcr6XQoG
H7QG9DekmPVwDbe6bY1wSUuEZ4ewr8SWQeqPw30qSmUOiFnAN0ZWC6MmACNNca42R/Ty6f2gK8yy
t3davYdPQwjcCkQjnqrUfbYz41zek8xqu/NAgYQVGniDsCuetGNMLim+rs5VUYqRq3QRfSUR3g0d
nvOCUK9/cCeuano490C/PQKh6kZQzOXiSgHPJQT57/MvxEKDM1AmAByxUeCm3m3XChsEdoAiSoq8
A3eO1gM2EmLl3yOaLxesTlVmtfsmNQOxsLED5y0Fe8yUZ6EsCofbVcG73iiKfsqTsKW++ykCo+5H
LatYa0HQiU2s9g774rryoytQuq09tPyYsPgfRByFksuTWeK+v6YMkxCbbReE3gmQ4MY/CY4t/+r9
SRTQT22zyVJTTj6YGInf1zTWxfYvk4pz/Hc3S6EQhO/EaCbGlEAqJiyWMQbCLULNndbROPwtl7Nr
I7rqiI8FmCzlcFitVR5H+lHUJtWS+1glqqijM9d8MwTdW+NRlOEKt/MDVFM1bJf8+svBMAuDACCD
BnWH07ceJJEZI3vIk6O723t0JXYVgJDa4Fq9xllly0Qf6JwuUQFb3+9YkJtHrrFvj4BiimOja95r
mb5zH/7TtqR9SmLujCbC0gtMQPJjzgq+/oZqFfhmjZ8pgnFmVOCVN6lrRKxqJ60SeN0XQZF+pePN
V5ZSK2p7XEw9spiduUjOkDaTRfyvRE4cvyVA3R05bmtdXj/plYJuaM3s7ZjBQcKrHI5FxrfwSB5e
S7abb4b3fW9P2OoQW+z4Cfn3qrgdFUI6VHkQpipGao37fqh5h3l+xpC6ZR+/Q68kEDquhZwc7PPJ
wc/3tNPYqrGTKN8Nx3Z/xGvRQeD748iJJAHHU54nrcSbE/+WUyp+iMwLI0zetrSZeG3zIAAoFkhr
2KUL3JrPJKeIk7hDhARCOs2InCpOuDJNf8JuR+Oi6Qez4LZw0HweyEm0B5PvOp457lNFnK2GDfeY
TvLvef0g4UpgRwqmLBS/diApphKpdySLPo0pYAEnrO6ic6jkQ8ndIAeLFIYN4xcSlUHQM9Medfbv
0KLahxX/hUJJZ9buvpmo84pkGLhy6v+hXjzj83MBBIrjUdGzTB/aa+9Zzwc6FL9+cSdtfCT9ER0x
eRBe/GS8P4OKoD8E8KrINO4cHuBb7Z5ODAJHshUvT6jBJhErcT+vNTAfXpxtdg63d75cr9uF5Vij
HOj02JAnOpttM8oNJq8NKBTQy2gpU3WvZyEq9Qgxrhhvmqrg8fxvS1RLDNqrfl+4YxJulKqdcADp
gm5HT35wm9IjHQVoiTZtr5WIfrgp73H0qDUu96HkU8jE4srLds6TS/vl8uHnMOhQwRuxtGghhjV3
SXobOKTi/EH+i3EBYNAeZToqzkIY9vVCv/tbj50mdREtiCOG7I5xcLsDRdlwmh2bcBeenqe4xmMb
uj/sqrODt5QSMutyqhenp6PiXRYxo2tWVfyOr2v0bmkPAullJeAStB7Wk+Iw8edioCDeN8ZoEhzk
C0VjrsVj5A4H+VSCFkwe2bIm/Ob8QDysJDq4Qf+L0kaNtTfWsCnGFrUTw6Wfc9oqzj7EnOGo9cFG
l8MyBifJr4VfYMmh+2U3SjJrz5afDPSAOYd8HkiLj8NM/tYwvSxHokx/+SsrShbZKK1BBhfk/rw8
X1i3s8nS/W9bv8Pz3U5aihM2NFw9qjbA3PdLJIYiKafNClUgeVioylqy7arGwALgajCaTr8D1+NA
OPCNRupYEBOJ8JN1c2LuOlwNr/JWOtETJv088mfSdKBDitJdRZmnPUFmk3O5e6+ol+tIX61hotbt
7f4gb/oxS3HC0nickM49C3wEVGC4kI+Yu0tI2PIjfgzpuzr3chOx8r4upiWNrFtnwKIdVLhzZ0km
GIn4SKISw9TfFrus2JgyMWbtrkn8lqO4HOGBat8hzeO9Z78e5LSLdTH/qXHSVOlILeSapPpNa5QK
TrYRt8p5VXg+gc4ApBp3s/S/c1EYMrG8HrFKC82WQztLJbopGyX4+tNdIDHuIB+0IlZ98ECp831S
+4e7h6uGOWbqUle+KvzNgOUy1vphyrKkWQXVBLCp3/A020kPWv0G1tKhA6l820OFX9r2AeRzkx4q
pf91JR375nUDKahTX5A8Gjupm4wsTLd6Hz6/SXFjR8tmreX1u2z4Q5zn5NgyPjfNsI2dCPoov+qK
ij7ZFXFUql5nss3IC2ZUVN57uyi4EnMM4zlJBov2o4c0XRfn1f5VKRbTZTauC58Il/7UPMk/4fRr
Gaik1/pjrrLR5iXZnb2mfkxef4piGfDXG9sOf7jjlsi4E29YE3C4v+n/qo1/BZUkkJ/aqQAfzc49
grw5MXKqld3v0CAwp5kyMTFHaPV42ERFoi86bXjIMicNCD9xJWR9686ItZ4Ew/I8EIkcRl6hS8A3
AFgEl+fn5WvMHl810P68ZY+kkgLeNVdiRGsiYpuPfE9SYuU5erXudrF8yP8MyMFJ1bsWGjdYCmcv
W7WLuURuoUzaB8Bexm2g1FOUK6XiSb5Bd9LfDoVESwaCBU3jsxqVETYLPIFJEkfHeDFMDhrOJycm
WAQJF4yv4JUeNzTROs8Bg2iGuyhcGXC0KJXBiUzos/RCph9kVs1zkCzmWvc69ZGC3nzy4uiwoY77
OW5oRGg9ce4yWriLPjkDNJx7vurBQ8ZeyDZA4rGqHtPBuXwwAjRacreiD/sAacdBNrpcdt3quCxR
KN9OGWlgsxy5nwXJMNJBNvVLD7hkiqsE92DshPUq534Sq2shsYgRjszNndbsIu82DCQltLsGeFAp
p4kipdHZg5N2hXyPK1laRkBwNAwlOW+lZq5G7AOxhH56MxAc2Vw4iPvrbMYM+lHEXjvvJDTYTcD/
4gS3QHqRxK2JCVTgLCmaPbBWSb4ayO00IvHy0lyYWSzoRb1zxwLLHNJzeZzWoVEwmrqxyUkopZfX
RS7FvEIs3A+vq+h4P+1KsFLRVXDiA9OuZ8cuSimTY6C2OmteM5W6g6upCLpdZ6oYdEiWjTbYplkd
Xj+LgZKg5xT0lw8Affrpyrk3wIxXaFUO+abUl7muF5A/DJI7OWXNsmAfrznazl+FAC4OnaNiNOsd
36uIB2UePwejU01uiiunWiSbZypY96oAjGQQ1P26Se631NXmjYWg3n77DGtDvywGESJKe4EUhJmE
SEuKXpPY/f/Cn02ZdPAkpXMmjDvRvsBWSwT4ZwBh+Q2GkxUIR8R5gkLE+BhUInbE0CAK7/llFp4B
SPLMK78XIJtZVIP2EBYT7ym9yi+qhdvHqmXUjx1k2/h2ar6DZDdrxsuBtFN1p/M3M+t2OUG3014O
NNE6hzrzVpsWDsP5uNEStc5bD8F6T7AXVXXdWcGgfDWHv0gckVKn+y26+QVkJG4WbrFAOQAK+gXA
O3ikFDMujYt9GvUV3IVyX4UgrW9sUr0n0RuVW0TvHVjfxLy/DUBiLeG99bagv1OTjJ97mz6DiDJk
X9n585L4sqMyPRMVzaEg6O0RRRtTRz0aH+FF2iD4Kl5hgWBcZRtoiNbKQACS14FpSShqVPtHoDxo
EJIbd9yZSk+x7F1DvK7KnroQsehQCW713RMvyPtbe/W5lJSWKrHHYtmv03FLQ/NEbrJeJU247sjj
1xC322IyKjriMaiiizqUII8TBY55aenl1SI76DzixdjQIKExv4gHCtO8PjwU9HLz8HyIqShGgQ55
WYD2lc1VyIw+yfLqBKI4GvKcPD9WPGOkGWzKB5wvznZIzMhLkat2z5eU1XWPGwFdMXkLxMiKZ1K5
EufRkyIu1mB3OX9jk3oEpKLcbNWXU8sYiow2xb2c84TKJaopDGeky3GPwZ74H4wNpnB38OX0PycP
KbMktGwM1atzEYfrpio/RPNUv9C7P2pQ9gUtGj/AgQh4dCb+fRlBST0t58NuNRT8w5HTGlcBuCeW
sGN98K45QBfAzEAhszCBFtjSbvzX1NbLmF0g2DZtP+uYwEtReOF8kD2vYFWjdWVNxrsRGKLazfDg
r5KH2w0zRtUr2lAKkWMz//NfMrxxKV1okOyHxxBC+mTqxf4+G95sTZOvaYrc7ZbnT40ftNt8uF+E
bTx/0B2RAfC/xGSsNTAB7Egu/6ztygUijKObwGdzO02CWVVOwhC7/ikXCSzmovVLqP9WGGP7GLkT
ateI87YKifv0xDOEy0UGQOZhQt8WrT6K+dMQQH9ZW2bs+QEot973wfBVqzyp9Tt06woBk9TwrdX1
nyLwIKC59g1oqOfNrZquuDKthzvx0FuojCRZKyjobA+VV86HsIIK+kU69OljUxRfti9woLdxP9Cq
kVJs3CAALuR9xVth3eACO8oKqtzmTI+8khfW84TSj3+G48mm0Lq5WOS/0ESEf+HqfwnCfPVSV6Jo
KWri1hX/MfjnaQwg7JxghXlJtzcDrDWdNcCImSr1nyfnTl/kGse/6v/GsOdqC5kMnsp6cYZLTrR9
VWyYCNhOaBV/AX8Bb44IT0qfU50PqR5k54YEltvCQ8y2F3xpb/gZ7IEKe4mg3beExcd3kZUSF3XA
roPi+Xu+F0x3nnfJ1zszI2uYjaLkYPL7xobgWhXDp/HQAHAlYbhDt5jQ/eX/zuKN5lkCmT8GkVQR
DMlLNQIVYQ9QLr9NZifA4DuNk43uraumILvRjtGMjKgqCtmNqUj5TOYvQNDTCVw47qxFy7Jnu5QA
qlgySkVJU/r2yKMpooUSIaWk/wceFdrPPTKIGIcbGQwXL/wINogPZpvBlvkUaFAhV/kfc2r0rOcD
tl5ieKDrrqgmQcfTcCsWjJHPoSqgDoxNX9lRVrPXCzcN4K/gOzuDBG0UbpUJiLIKxcUV/ojqRLvr
SMT80vHqyatqkuyCqIwsJI4Y643JE23xmtV6Um7EDbYs8ElVE5A2HGusgRjhQsTn8hrxBa9uIMVL
7xYBRDZcz6bSHbNb/0cV9pr3/pjxygVnE6x/OwAap7S7HC8NUO9kcg3ZF8dj1omodc4x/V+KRg4N
jIRGW0xCXtXSfz4mBeSDElPHnt14l6YENVgvp54LLeonzViMarCCT54sYdACQMb7U52DEWs29way
AnqQDEropH9mqp/IBAbqn6Oq09lskZ8BKBIZGJEKBrTabNk47IUuthg7HG5i9Eu7vl8fmMy/nE4r
WOuuVtN7dgQ1NLNOV8ydkVOBTZE4iuynIDMobV1vfblQEwcg0fK3j9g9qraliYgv1fF0B1k2z0K8
PIxEOy1To5mhoLR/eB7U3AL7V6U49J3Xuhp6EvJmJUhirbU1bZYlsuMwAjjTZfDkNoVT1jz0JHfh
wtridG9afs/R0HmHHnDpkoVeP5ZZJAnT6kQB5gQfJn39MSY+vrj7DVbnWOeGspHT1oFE+Q/IxlAr
SUNnBt2E6577VT6h7tu15yIoFo0Z7tZwIDwpumFZwl9Y4Yybajdo7hfOo77LFzitMIy/e2ZoxO+o
4+YaiaQpkVU1Gi7K67uwjVxxZhSVnlfU3dXmHj4gex9fuMv+rp/RHbM4T9U+HfGNmTIYZ9uUIm0F
9yLAcMik2RXHg+5e9562U9/Cp0LbIXXx3JheqPZzZQgsp8I60+BJtSE1NyFiwRf/fgFHacPbXkp+
uat3WpxkrGic3dzOr/8cLtApq02HmVCyRxnR6ZbkVDljR3TKtvs2XnZEs0oUoQwPjglw7g3KIx6I
VZOe/1CPFsV6V8UYmrJttOJ3DuQnOV0ntEdzjdX42dMWDLNs2fGmLC170ECzTnu1rtfQ0kftgy+w
xGx3wJ+P9xJQVigXUd378vJ0mev4gKNEeo5nXzI871sUTcGgrt+bvj5VzbljC6JecmKwd+TPKMPR
EZrJC+YeAj6KFuURAKabcIZFPhCo44iPURLtWeezeL18CHl/Z72gl7SyPHY0o1BqbVBptFl3OvCC
rvcuJ0pvGss68fik899hGAre7yOlN3vI62V5nZS65IesgoFi/jBGn7OfaRtj+bxjgyauhwHhcF5A
pTrVbCZNKSSOZNdIufCvHShP7cJFEKu6iyfpz7aiaZ2SYrWLAmwBuPVeg42Gi+7JZ/jFzOEWl2GQ
DtChvN/ZGLYizYPkJKaHBA4gJYUrzJ5RqFBUA3AJddyR9MvyctSpHfjLOlioGNsDyZSs+UouEE0N
ezwdyX0EcURKFSufTGqyHZFazqpThUOwwU5hSXFm8fRLHP2movwGbMHet0uxoOYc3hYm5gbVN/Ua
fFzch4aQmhHoRwJVDGZU+HcVLpFUO4LtgE/z/LljBBW6chD/LZ+Z52tBJWzQnlHkDMaHg9W5ljtZ
E4fSEVLEBPtaI3xfiHeDcAIWGtph2nFO0E6nqYnbgaRUvzZUMcBemCZly/IWeOgisPHaQZTD6WHV
Z79icdWcVgus0+9farHfVtHRRTNu9inAh/WWTbue5gls3dub4+M1imj6ezBLJ0SK6f7ZsQiFt/VT
/Xu1bvubLpMzPL9/2apA2NC5Ye2fK+1Hq01vsCKGMlEEg0/5lGtf6n0Ncb1NjB/h+1cnNZ4/afy7
HbTqzqASXYiVa/iuArLgXRA3rH3HVLbhjtvdhpOgO3g4qSo1N4BwUTujF1MpwLrTf81bPKpLqIPY
8lQSa7oUafNrFFGgOByWxTvWMOCf8LeEBaKj8TLgshXznRfSfNSU4WdSicgQAvURrWbucLE6X/q4
x4B9gIzugtqNq1W9veUcCoDMSL+WoRaowTiwG1E6DdtxTJIJZlk+IxR1TsLGuDIiuo2d8nwg8vGl
FMWvocvqWzHlw+u53RWFFYblHZnA4RHFCwPDfEh0BbFi4BwGR5+lUrSTMqE5KeMufqWpXa5sUxAB
fiqR6eeehqVZepdPPhlQXeYdGt/g16UdLkJBV0wnbWbew6iEhbbHkTjSgLU48d+ss5P2KgK2yUi2
BVrKhYHBJqb3xu8oXBPqSMcPAKzZxPVQJAlvjctAW9+YsdqCPdOspNod4AXtYDzTFRrgET3NLZ5i
8mciMIF/iMLOJTyRNc0wkBnZGUDFgGQkIiTY1+U+1RPuqe4pDt+oK5gcy6lPL8pgANvLcakgUefs
II3DCyAfLK7OoeAklT6nWRJcX8B8GKBTY401G7XmQcZ+RtPLKfuWEpUluybkXIoLlMsmdoOD4yK1
wOhiCfRIiXH9Grjwwleg48UEPjFwofJWt9evb/mFniMdBbllpEATW2Xmhq7o6ws3tx0fiSTyzMJX
/qa2/0zEfbE36+k4fYMuPqHx2rFS8r6qlGTEXgccdKEE0QN46lWNzNY/B7f0JBAag/nDFn/CNU2w
7zWMVSuR9x/zxDKG4nGKKqsA2bECcJ//J4ojiPsXnCq99ijHHPHLR1IsZLFzBylOB+X4SHkUiuad
+EsThc3Bp5YecqUJdxaCLfjS03viqEYrUS4rwZVoGr/SdmhnsFfFCK6jH5rsDZgFmdTlgIqawaxq
AI0FgT463kNUX2+tlNV34hVLiB4jCCQuba0XvLzZgamHlBbvz6q3ptOETzpj9eEqHtgF3ixwNqAG
OgQGy5mts6TPFyHZvQWRSKMXNDnBfgKo/4oHyffECL8McHKfQ1jcUQcLduoUntJdSqhus97zVV7H
fFJ1uD2jYBLViGqWtDxWEEToZr+cXo18FrSl131MuLxcv7Iytj+YMAknxtndhYKW6RtTHMtAGz8J
I6ZYbcmnwQuNWS+3tr5IGpvQvcUNPTbyJSokjFAjuQtL5W6SxO9R5GYiWIGdHmhx0+PCNwmjadLx
muqFNQEaYPtu74KmSAB4nIeq6jLo8Vg7apQ+YTrE0GKL9TSbTKAjWNBwvFAwEiT2cTExTiCkqIOg
Y6GrImywL496WfHJYmArWv5fnliKR2LiP0wyyiqZN77nUk18kGqH6zvXcqOPDRHnrhIcrBjqBVab
NgFN3uq6Gc2HZQdE3Ita7Kn8OiFPwfCBYMP2DIA/9qToKxH10ah9Y2OAhfmdIEz8FjaTYXCTUeIv
x0UO0zI+TUWHT3Q/XYjemRUYQIx7KCi52r2w0bvsj8IXnwFO+Gg7+ailzInetDhC5RpeUfLp3Hzy
daStCX1+aID/cWhCA+I98GS1rMmr71kMFfYKOyfgoKLWN1wKUlu40vpaSivnGZLHUPN8+tJX7JxJ
brsKogE/hNfOXHXwqpSXK7eWWOw+h6vAgNaPeQvB3gqnp7rXGRV5uxboREy7JVhlzDSyII19J10u
s7mXCvK6/YCR9X+skk2oyuBhZguwTLVKgxrV9KFI/Y3mR9JH16Lkdn9AbTHBzaGy9hdpg+4RswcH
iAzT9WE4maI4PRdT22lT2sAMO0ykz3hN+Tqbnn3FkjQaqFf6MicAyfgalawXnTm7KThPhIL3GfZt
x8aS9q6M8a8WRSN9vHETW8Tu5see5SLXF7EYSkAAfCIGyoj4vm66UyE5zOrGhzMUoaiJ+c87DnRu
PA1edfEorQC21j0emoEjcvGmeFW8J/ycltaLr/nOPy+LmUZcmYYauHLSF5MaWQ2D46PTMCDhDhbD
5N9ZS42z2e8GmZCUCeWIWgmH5m1EVdNWZsmRaJQfCvx7wffBZ4OiEtdT+v8+bPrXs6mRR1ytjNQk
Ok0MSkPeUsqImq1OufkrRGPDa/4XTVFuVMWoqIywoSAr8yuS5xrnK7bHZpBnsDVlfnGiBNlNh9J/
oiRwmLAGe/pT4Vz6TJxLSEvLVZN5zaNCPRvMNYDUje/kavpZWg0Uy40QSdsiREMEnAvzIUU7MqQL
o8x5/5PE3fdo6rKKInR36/ebKl7rZEwye400MkmpbRFDpz+c/ImgLUFpd9dy3qyDQSLJOy+Hue2R
WIq6ex2cJ+0RcsQ8tIQxA3NaQnb32O0lHzyVlTsy57pdcB3TfI6E6xCvziIsUooRWbbb7VGfCAi5
ZwuI7POj5FhSjKcGcSCrdal1BRS1PbyJouk/idJl7Q+ShlTbbujcU/eoSTkxvhGWvO0HXBtTRz/J
KABb3GO0SIoLoLufWfrkmVKtnw1TiZMDaHBzQiySdyqXC3/k96jq/M8KHpTeybkr54jfUsPf0Ovw
y6As5+oVa/i+MsnMTawcMKx1tRxDPiY61nUp3tEhuVYdS0NvnfIXDo1sd4Al2+j0Uz00b4IF9Xqd
nT+vX1pAQLK+GgAzwqsB+uHOD1/HVxoLJK9bXuLt5R2OEAP3nr6GYvRfffHfY4icRr0dOHtWY4Ti
t94+I14RKWY81H81dhe+Camcf06wwR3TeLhK2JgHqQ5w3pWZCLMFuv1LiMyAjGrdemjbmM2h3KLR
g1gyFzfLMOC3LJZtmdPXWKBNSa7yLG5lpNtqNmOlGI8cKz0BdyZ1T/w12ZTFxjrZi6iyTHPBJZg1
Lek2c+MQO4jz0UHGSrIk8CVvZkSatiu/pQGheIZtsFuE3jzgejwIdtG2ESrT5K0/R3B464h7eVMA
TKAy9U6ekKmn+recS7H4/zmth5+G1iKl+6IZP5lierKuHmwobMutnrbxHUjXZ0H7t/juNWRwC20E
jgO2+mX3e7664QhXlFoQjSi872Oc7umnVlulnmSNKm4uxuyXhpEjhekVJdfWfXAa1H2vnZQxYl66
Qj6jew1TOLi3IMOYpKVO8dniwSpUVm6H1kY8Y6SJskFb8Mv/TqWD+xNIvcpKcOQejGdcpWK7Ak3/
gkt6AH5UdBYNZDVwXgwbm1cVIuJWATraXsabjuTKhR+O3Gbwt/jch2CAJtNvgDo6q18wRZ2zTlhw
QT9wV1VPvomjPSULFbsldZ4/Yak077KhbFDzHzthTVsjQy7MRcQtPuyTX+adZFnreJi8KOSqHB0L
Yv0eHiYa+MUECChWNlNKhJw52ofDeZEz84IvWsMcp9Wrq3k+N+HZhgcEF/rWy5a80YHb0mIgmmUS
eelQQh37fHTcpoGIegTKxLCyNR7hrs9toEihHS0Uu3uiJH+rWWTOoRFj9/cScVFoC1BgY2xsx1yL
r4drpA8rBUPsiWfdfVsjFWl0sRWqAST3ug7KEj8p4BUdHLLQh5L5/w7HLx8uDPLNpK3nikrAzba0
2FdipiUKv8wal0/SJrP98ZUty1dt1ArSkZlAhAL0sMTXWdOg5XQxiB7GAbVN4SaYXXHNwON1jmj4
Yt08GMIltoVHEg1r8NRDVN7+MW1L3YMffAv2s8oWoxNbXpCR11M6JprLx6G7s/KP1ymEiBN3aJz1
fknUDEr7LNbsYdrGuB7Uvo/5AjhmwFG6xJ4Z8UuAawgnFHRjqltG0oBkH0gCgd8AH3V6tKYNEEce
rr8SSChG4J800TIHoM8pGtCAQQiP+FLRSM8Z8lh8X4xOv5YVXYMPIGhC22ZVKmxouIfkYBgbv6F5
dmQuXnYG/JfpLr+nMEo41tY2xq4ihV3PsFENi/IGFtoDGAMGgx+GF12NzJDigb4McmezhXZSuqww
MtQ48c2ZKVLraPQKObzmK/VK1wgN6XQC32ZV/uJLfdtzcNryFzpH8v9+QckcH5DPfhOGVbmIGH58
sfYm+Z5Pf0Q+pWSG8gVbNOrWoOSWtR10RNYiKYfgiZqgakRgUvtf4KSVdr83aUP3oafv4biC3ll5
TXVWl+p8FtJhhBkL8i8ZjQMKQv4UjIqSTKw/X5TJrSvOhXW7QCatueRvyt58PDSewZCIBHjJIHWK
Q473MiZE/b6M8PFAT/NeAGW3DZd8yKO63J6MWlYTtlRrnBC+WbdfCykhfSNfRJHnUxnL6iy1Somp
ZqFGPj/dLMmxzH8CKJ/+l8UtYbZcquN58Sa1XCDEbFpHSVZCuR1naq085edZfRGo1urb71AuXgpz
U6FA2bUQsmEl/JnoXO4OQHhBJT+AClvY3eWHm/znNxKxwHk7anLiMcE+SlxsC4T7K3rySaPBUnkA
a0Kext2fyMq1oN5ww+KIHFRQ/iK0+VTvIyHdZEMes/51PdODWG7q8Az7QFdgsvD0KwYSH4OYDPKz
0/v2J88hst8ItBWocmn4VyNPSdmU5RRFEKfH1tLy9bdDgawce/MRFIz127UegWMCMsF/7R1iULyh
QJiccTql0lVaeCmDtVoNWYCYnKZht3+yWSeHgkBzewLaDKWvFKB6247ln0y4EXduBp+mGtZ5owzD
JmcVnKXBinxiUIOP4VTLWoEzOlRK5PPZmcOfXkD/EDtxGT7Dp+0dfILGi0cRBZ+nj9rt7Wr3xey2
8ZT61lX1jST0Gt/26SEvXpoJbUw9Rg6Y6ipoXLtf/DN/VmKo/rcpuKRSJ1Wolifno6QOr5YyNcGR
zWvSPUf9k30spvm7PQDdwaArZcgB1vmp3wZkaAlvNcIZcTDLvIsMkLDGwzgH36fF25SIq2/SiLBD
g1Jk4SgVMWh2Hv6Y4cVmbonlIC56WuSUTadKH8a82kGBN4TF7fFNZhFotm+qGmXPuGodAeyZClZ7
l9gK9FY8eMls7oBxeTiGZoUn9LFrt8Ex1N5Bt5iEfSOTFAyLHwYQBj5vkr9zYOxRd2jjv2eTgzPS
BjghnvDOPF/VdNyxAbZWdkPUSsUtdil8XScj76O2XbNU5WEHK8aMLJRhmDNcz/nQ4xmwOGkXf+7A
/JoXtNijZarsgRLrbtK84Wo/qx4kMg7EnA8SYQPkSA7c3msd1/pBUQ00xjy8P7O16pClq61m4FBi
J4uFsquosnCyylJBELx7QP0t65xx30HK4rXuULh4EUQBM63io45N5f6goJKl6RDOvbIvIz0/bmRl
A3kGGZcWOHFnKbT8eHXQPAza8R1lOS3KP68Nv0jK61mew4wNXBRsVgDN4KL+OzVxxqBBmbo0XsSE
ASmUepF57XUwo7hZPz58cmrMKtDH7xHiswyqqXY13MNTpMfEkAzYkK9MMyTgjXZPMsSX6XkVWHky
Amltkt182YJm+4NPTLVEp5OXZJBYWXdbJm6S/BnDZT9Y8FpiA0Gfsoc4JHR8RAag6MdTiqdJNuyq
HI51RRvXvJ+h+8GJZnd93DiYZPaAps6XR4JK6CatSOk65gPFUF1bwJlWVpqrZnU1sOO+D68GEP9t
Bij6Cz9VgWwy1JQITTFbQxg3oV5oiWDArtTbzLk0eRahyfMsHV0S7FWzFJPClKoa1/486nrvyh9O
6tNnO8Le11+GKm3R8syb8cM1yBEHjq3q5rY3x8fFxE3DRhgsFOcGZ0DNWfGAmMc5jopfct8zM9rc
l8XG1ghR1KfQ6K4c1Go76fJC6ECoHtbu+qCDk9BkLw2+KHxK4UYFVlJyxRpr7WrQM8BWHNz+TIvs
6Tai0ZeTI4VYr+CJV0lFw8ZQGiDA0lZlLAGE6B/R/swzSkMNB3z/KZD9rs6l7Iv7DJj2WqUT9Mtk
msdaD2vn2j3DiVpLLez8YMSsFW3g3pnYbG85myy8OfabbZrlwPmz0eI3YToqjnCHY3Y6eT0pYW/G
11QROc/0C39sc0n/IwUB2vmDzyXvB78vmgNbEFxiNnr7wEaQUDDBH4obQU8wfyz+9KGpjbUEt+xF
HCla/dyj2Wy2Vw+J3/lPoiy/+k9q1fdnR9T22goBzE47GfSy6HNM1f3jvzVBeZLjgM1PQMJV66ty
bK8Gf3BCNTY7sriTrLQHcwiwgLHAOgCYLouv2uPw1cDKjbMiIjMQg3hC5ms1yWdV0D+DOI8w2mgJ
Rx3aODA/5JBVRbgNG9/UPIOtxMQl5qCkKjOYuJHv8dGMSV8Fx6YWlpYmjerIFSyN0brX691MfKvv
2AdnPZf+HhbdouqNjoxOf92Nio5d6f+8+zTxLzlF/+T6a1R8IQKN8CIeZsd3po1Jhg2SLBkZesVn
/hi8x51nbCB4+e6pFAfNMJQjr7qejt9BdRkfWYCXGFA1QijwLoWs3peaxqb4sp3GYXm0XCS/GcSE
dnHQjx980paR6kwaaHDcY4X+ioXrD1nsbK/STLOyzYUk03jYO+n0o91hTWwUki2iU+BN87N49koN
u3FbssPCfK8ipmoq3BEm6FUUG0eBMu4jlqaYByO86mwqFLWkmGLdBQEYmBO/O1xOk4KkUEIMSMQ9
ov6HYPaMAY1OGsDAK3jJkaOJ8uMJbAYcSTeMdiGAVNhK4QK8aAHbMd4nXwLeWol5zCr2ESdODqJP
ZYeXJYIFqmLJR/R2SFRtrlYNEndj2eK5mgfqdrgBcU1YGXXeX48OJhQSZo6+s38z7y/ma0fms3EW
yQPQt9KvVohon6/odEXzWQ7OOqEzDVqwt3yAzwlsa4t//mrEjLX8MK8ur6NYWurl0aLwsuT70ic1
MFMojkX15Hery5GNuFtWATluBDOxtjPJ8AtvdJm9khAnUVr8cNjojLcbzDUm5ZpTdy6noEs5a5tf
YC8JeHifrCEFSUAtMY3sg6oePoVymCXpSmXucEyTazqPlZiggxJQ0H+k1dltSfJ+jHw3R0sh0bed
tuETS4AgCye2IlN3vl9v4pHEmBkk7s4W+j+xei/srWKuOBKrI7GMgAfV9p5DRXE41hbLU1j+FC4q
jKiqdHugcsn9jsKty2z5n/lJyDxfelojbHgNQqkOHtVD3H9uCv8kuq7gCSkNLuvUQndR8hGIwzET
v/pMWEDdXLGvLa1RHOa4urUEfry42uOMJKJPGXjMJQr7rJdYGkGKwFcb/2jrMjU9jopgkVj3o9Z/
/fALFuc+x4iO6nKiyQV35/cyBbKbjdzYndcOrjFwYiGvH85luxW/KEeZ2JhzFogfv6hH47wVomtF
NKhQnxXjrcrw/PnnJ4HyXvUILwHIIe3aK76lyh1/8PUVOIIWB48Cdo8dAVcdwnbheV2FSJnkjhGQ
RdGGy4aDgV8In5N+Rxkh4yDuunYLGD5rTjmLZRknDdHdUEbU88thfNVfNGaQC4a2FUMeVOg9MGU6
npTJxbZBhVVc1Vo6Zg0ABG+rJ+VjKvBEZgWH6TEZUePzx4YL4HTDWlaiVDsGYEPcOyMZlWlJFQuw
NeNnBS1J2HwsjnfeLNmNkhXcdHQif3kmGZwG4f5jUxkzHdnw7vOGiV6uChWEmL4gc0JfuyNXQH9U
goRNjSB68+Ew/Bnm5Nw0Iq7kctAl3DF/X5dUQaJDLSRtirH6OJkVCW/xD91Iudcn8LIRjDvSbauf
AVAld2k4CDtVGgLSfkGwrkcDqVBGEKxpze/HtX4F+0K4+7mwnQIvOSUjb2lLtQqtAqeKXLL+tNNp
fwauUqj+z/rybeoiaPo+h5qxqTIFVtDR3AymdhyBEz7FfYOcX2JsWq9NLqNR+e6RvA4slPXJQreK
EprKe/DyFQ7agiG+4kwVKehZwescBOz2Yo72JVcztzHJN9yDUT1nEGnltOA+QDBmKLu0ukvaCXbf
4CDuY8AW9Kqo5kgb/zz+mZRDnQPx+HiLMdAd68bNKqlCE14qD9M+yoBD//VhgDvWyvUG9JQN0YbU
249kemoIqLSLyMeDOkkrA0jKgIO/QhrR0xPrCJbbM2zqHaZvoABaiyM4N8S8Dm0PPLv8IG06iCTK
bIJcv0uF6p8sGJPWJCtV9qwwGCNI2XOWg0J3++cll0lAfGMbCaxNtbNJeUk0MTSVIjL0zthmOWF9
U/M6BtWFgiO/WQRHFkY9HS0ZWPUcOOuiMzLb7vFTvqGS2olQ6XkEAg0lAvFrwlHd7Sqqls2QOcF9
hr2EToUIkQzSlMOUGN4FFdM7sge3+CKxHkJznLIGkdE/voHTORQ/i5R6nZG2eegZQgx3+nNiSRg9
39/QboKcc7Ar/PcNVsYyjxwPrHdfezw5aDHYHtyUq+db7Z2pq7FsWeNd0uzypZoIXXku3LngmsWy
X8YvYF5HobOdlqIoCnmoKhn7e0yIXW63scO6CW4Dq/0JfYesWWletB12Qv6fEip9n31Bjen651ec
fKKuj565rtwN1gxPy1zfqWzUYtC4dWcfaXOrlU2lnml0lGvtMYoh8rbD/RxT6//46w9DnLK8Nyju
81QpVTVr7Egbw/jadup2IMw2rXxOA4eWZtbNrJWnY/tkxcZDX6O66v+WeIdRc9sFrHpxNPU+cYGH
zp35L+l8ceZbzwUrv60MJnCk4owRK7cag1iBiU14kw/PsxnrCMgVD4tLvlVe0qc/S32I9NpggaIm
TJkfKqzZsPXOIicibCC0WaATUX/c9a66EyRiyhARyP4evYsZ2W0sBzJ3zMqfZfmQ28wM4/8VT215
gUcqda1z73SvR4b4TKtsCiVTcoL1CyYor+5VPzdqabgBMEgqQAq/mmv8OWF9JbEFU6pOdngvQKeQ
x2erGGBkVF4IU4SP5Sd9qzimR5SsVbV4Cr/dOkUhvDd1RYivypslx9CM5lEMJHIFNE55+LjCMocS
vIWVxhLS0adwZxVcWR6xzSf/KdH/K7h1kA5el/kzyLW1bVND7XAq15nxLkU5vHt6PMHIIYVEq4sB
KzuJOfcPvD2skytq3N6pjccB46oVEFGeyKDllKiG4/2cNLISf0+s7tDTxDQ8bxCCwFKRRMqCImTl
BA7P+KphmcC/A1HeMrRt6sVlRuOm6zb2Hcl0+xB8iBbuMR2ltkO+1s2yiBzmB9GVxQlCj8GFQQp1
ilmbEOTe01VyiHDNz+w0C6I9tU2IQIxHEyGOykxAPH612Dazc6TF0ukdSZ+I9J/GrKh9x1Z5sHyt
V3SW0dq8iB4o8kzdLZ+NhqGTbYlmRN2YXnXV2sfyV+TMB+qek2xhygg6ZohsqnHDfqbPqqVfHf4S
Jn4aKX1PMZ6N4x/K9bHwCObcHhzgZiNuMViCrSUvCazmgqzi1cEX3V24aXvs4t1QsIwN6juLiMqs
sE6mRljGHm1ze6NbQ+TBIklQoA49C4Wt15sKYU5aoAiZQPgaYMxBxnaEY8gRNWW98GH8H6IlBsA1
Abj+HwBRJHivtxoRo0TBc9WshRqWnPTbvDn/5HnvxRNKaJAvL2vcOoT5+EVfKBN/PlVe5KRyzGIz
xE94rNLX2UFdYQuExAx0PIUXm5mW2L2u9LxLgIZHEX36lhtgQ3dox5wMizjbGpghdMLRrWhQboVe
TPRb7HcjyePPd1GQDdC5tFN41UkvZ0NUmedktCZy4aww3qJNEQ/ES05Kwk+8K2x/AjMtDmzsI+XZ
SGLvjuMkMzH5yfvkj5384x5rwG1EZcz0vAuTXZNZFKTj5UF+39+SYhJeWnfxnXMuWz7mCodm5dQo
s+Go6jnCfx0sK8YN2VmkynfSqFRq3PJ/zrALxlLsoC98E5y3mim7uSOeOuLM2oEsi4I9OhpgtBXE
i9PUE00fLGM9xJyrTkeWuOjrsjoI7vRFYuBwGYGfdh47iEdlFt9vbBOzn/FN5mlYUgwCzMXQaUqT
jfw8YhLuJ9SQM6RnUTRX5nzk7+h8UH4ExB2s7//k0InDfvSILGjhxBlJoZxL36Dx1Np+RBi9lHSp
tS8QSdicD0Xp2QNgqXPwVnaZuxD7n6+Oe0s4Rak99gWLsaOMqBJBeZtKsQG19KeVmwAF099Axr6g
sVTappGHUGfFZlAyLHub6RbAogPu+I4YPzYkeYQZsq0u0GBKYhswZdhLLqdtZlw6fjKjGab7+arK
HsREBXCbajx1DmdguI6B0w3IQJYui2Nww7lMv8cuveldvbDU2hh7yTuYsKF03Z3O0ekt3L9EGQ7p
XAfMJo8FIIxXNhZjHIcJrwf9U3O6qtuZyjqYzbQCQLb3NfsZSBWhiHilrg9TUehFLdPkw8CGbL7M
Bgzn8E0MIBzvJLmTW69FfQ4aTYu34vTu3zea6YA/Kma0dU3sunZmRIoj5tfoXVXPXvtaPmsd/vqd
+ReHSbYK01byBUV1G+VsHTbtLE9VveBRr+7kTtMFrdWBjgJf8WjT4Pidgu672Nq6wuSLQrTfX1ju
Trd9FjozEchIqxSU7vFWSn5Xv16V074yNbvg6xF5H4/d5448V910Byxlr9WB67kA81LUQUKUmjOT
U/Q9liGji37TVtHwy2VRRTO+YTshPyLFFTEVDvd1T38zc6hwt5FvAygq8fhcvjqkjm7IkN6lWi7P
XISPZju3mC3VY4VkEwKv8RP4tHAKabUGY4hhe2/WhvZyPccyJQnuThbL1STXe3nugKPPYrYnJVds
sy0uiGN6LEiNW8wTFdz+5rho2fvFzkkpUlAY9bo/kBMS/xjR70Im3Y5ms9tB9Q3WLl0qyniaBw6o
bC4x2tH+rO+hcq4rjUBQTbwJHIOrvTihkKi6GEg0U46i0SYNLGH6uhlbmpyImZUROIiKiym39CWj
Zuh1lAWWQGBrPvba/j5z+EJKz0ErebwZDIhAUYt8439aup/H+gT/OjgI6aVym8Kv1L9WU5Xf1RXv
J4eWAZgqtLIwwwSGeeQQavCbRJQ0TxIPo+eUlj7Szs+WnxrGfWsKf6dO5ibwr/P1LrGb8lwlFHLL
Do5vePufSWHXp1YiCzId3SjOTBSwk/y5lYXanUUcC58MEaOeq6lxxo6vMON/EUM/ao/D6J+nPRqp
zzIV7L3YKGgMglxJQX7Q1cpMQ5zHIajGShdahs4cMLaXyZd+uYoWkg/fu2jemQE/nsPRn0ypW5av
lFLD+zit+OECc6jHGa8XZqgGRtDgOg8iDTM7qZgeRaWbdvJjaGKmD6eTfuB7oOVGSMO8kNBdbNGz
QKUYzd4/9RwUxqdaHKhtDmxayHqgOLno9HAJUDbcSagF53qIoNsOZyDcZbho55kFqNLBlsHHiuWa
dOnGLRdE2P6Wdr9WBsZoES+Z5DvPb62sCDnrwRzn6LZkrNqKubk+V4IPeCTXhmecOah07pOMIYf7
Xt/Jn5PEVpFTHBo/ewmEli9tlFyGSP3lUUT0JFwHpBU0xB4EiMTyHIM42qw7wXZU7Qbee+ZgppyC
0xar42+UaJzPDPolbYfjFp/LkUmazI9vIUyBjIVVA4x6mztpCWIHDYI6LZkZwnhnvWIhPmdf/vYd
a24NiNSdW3vrdANp8bE9XBWmwkItcR2M/zAllqve9OaCpuL3XBYWEve+pHgPNcejLN3lBNkXI27b
xZJstZghmsGv5Ur8wxIowZjPCWDDBEsMdnM9w2X8TJTXGajdqC1eeyTCXYmVR3BCjjgV+t52NxRu
nz6ZRLBsTMeX0LQjuqzWxPzNYDvSZzDR0Nvx0x8Q8J477TFMxDwytGpBo1X9V+u1eQAfLEuyDvW3
CeB+0SJyzGxhdIjsrFrR4XgpAdJc703KBqOYjh1PuNOrtwUYM/AT9DKpc7f4DpeVyy9TQ09Hrz/d
rgVNO372Akwcdsgq9SFpzDtCw6+ZSP/HH73XQMDQtDVoQME9VgQU5QbX8FpZLQHtqurltHJp6ckh
FXlp3RFv/+5JiCN7XFbFa47mbpIOsz087ksF0qOsdwAjcWdaxJmtME1Dmqtwg0keBHcSaBxKAvOh
AzE3mKIg2Nr3AWRMjDh72B//dB3Dy1fsa3X/l87+mIBncLMEPaF7ZxqzUCJaqgvIoaCqNOn2Z6fk
BsX25CBNR5gtx4dPdgnRBCmpDJ+I2EPmN4s/Ta0aMZ/OVSGPoltkdz0Xm5dkNR9/kcsGEjkaWN+w
b+w7ZNAQRJ/0Ewi3G5ey90uTDRBJ8RSeUZVuA866tv7IOJ5latCEFQRhblqkLCQWnHt39FDXE7QU
vj1ncHHkB8R5/buIv3Q9fEHv8rSCNH7RyaqkO3v3C+LDe7HhnNFbsekhgYYz7OvtHi9qNknry+E0
wXYRkmE/wj3Ths27NWi/heUedOaSnSue8TjPwHuaESkMjUoSCEnTbwQE3PLNCk93Lj5oV4edJ2i7
mswTkcf/9qA2IpxLR3muxFrju8hZsT515XZDIHM6lr8sYPXd1B8Sr351w7hB8nVlOMkL928u5ipT
1oT42Iasj03dk0CyNIpKzb7PpdnX/p/NuC6VxJ2D9Og743uLeqNfzofswDZjGEYA9WE+fKLgVnBM
9vnIOo5CGt+h5kuAobZCNvEKlmjcJp0v5T++rNJTDZNhpAEojhTotUc5dIqehvno9DO1ZZMLm0yD
yZBdf/2UxgFpxh4eySMWDf1aMSY4XoH3Gakbu4JwxhIDxv6EhKSTCLjrgkpnBA3D7XzEzMAbbHHu
wWOBIQxbEQfSzqRQrIEG9UV4VD3F/vdeR3u34A+3+xXm/TlrlGhg5FfA5b1yr5U6m6K+KEuZkEYY
E2awI4QmwBac06Ddx6GgJtwdFCHaaODSF9mT/oSbeOJKwrD8axZw4FxK5AYsK6qcXGIJ1kwi+g77
8bBjC6Rc54BpmjXvspJWqYldKx6bcKJHzAFSxQByCDDrQyKGxv/6rNftbVdSd7rKsa9cE8VS/XOk
W234BFiB6P8LbiHInpwi0jDmptGvbMfJMkx0HWKm6D+ShXNXtuA61Y8bkM6Mv0Byw+GwcwgC/gzq
B2ltKxicyEH6vwqYDlMOU/SkqR9Ze79pYTkNqwkOEFQN/IvR8H0sL7s36/yGzSi8zevkYig4Y8/O
yseXR8n58soEk+bMpxYBVj/LTez1kQX3N69Pz021stK6/r4VpdKwFvJkxrGNfL5JJMZFoMHZwJnt
IDBHbccxrYTOFaNwwU32IFYUDmEHCZegPKj9qpppDlFpp2ghDszuTMVaVZpInaY6+kNF0b7/jVpj
ui3xjihPX/5B8RN4wQdjP8nbr2rj2KG2v9WHxGpEFzFQpvQh8DpUoRuVxJCB2pTWalGdx26k7l7k
2tAsr0MSxCZh5HWqCNdCMZVbG0Z9kICqNTBBsoq91Yq+MWfIEslbeBA025GE4iR2VS2Ec4PuPgYG
jUIZ/Mg/JJxdhjfSvEgN6Q2xs0O8TWqJ+W7C1Gf1kgRyk3PJWpPGIMDceviySqyZRYHFutUx4K1o
r8eEpvjwTJUep0WGQt5vnULGg2cj6NGyaLRkyDmIsYYPiYXEy6qx5u6TtQ9uiI17+zVBh/MW3V16
k8H9aC6pYE5F8EfsX88b2ic09itIvzWWtz4NV6WS0WQR5+JG+lBCk1dc45eur0WHAhgtD9TY5ZQX
+MkoktqNtx27/yakAtoZOKUvkXmS4csz1R9OnQFOsrfgqoTseRgB+AUC/NG7Oc2D0AuLbY26o709
p9EKbntf/aibxC4/WBYs1FmB0z12ZfiKqKl22gKtfz1dirt+OBy3udt8gPiWlZh19STdzQ5DPECO
PaBijJtgLBNIrjxpiFMt24qCvPaGe6XmiEBz0c87nEb5UDMUi4zT+bBSGOOTaFwdsEHG14Mm9MeS
WSnDuP+t7YqBTZB4cTi83YrZBsUCpYuhG8ZloMf0MIdWHsGPijO0F6810GPEesdU0iKRKU+9WHn5
xnAUTbR39RMWFdSbmvVQHf2k7d5lBv8BDS+kg7P+y8aPCd1jDu4J8FPxImRr6fjSoz8Q7DEvtHfc
ghChHgnm6grKqL2lknqvY3w1lc2c+lugaX8Jc6hZPQsqWQSiyUn76aWKS+RbgiY5yh75X03DLe+H
lrGehyPexkf50aOOtnk8rDMjZvfRQ8Q6nlKMd87fhLacVEMj0r4tN2T1GKYyR6h2fvNx5ItIShBj
80syeZeCNjC6Bi3zMPkjzKTBxZgiPXmp30fNd6Ny1kBx4MOtj7ewDUxUWcewQ7mmGnPfX8KO5lbz
QH3K2k3qX86ZRMuyw6x2eshINxEnvAE0owVwlbeKB+s5jcrJMx0djVHu25b4JkZTVgNhc4D5ikDL
Gh4T4kWdlvU8qxdBiZM7yc8kqB8Al1kbfNVR9Pkl8LT4iSKWzGIoDTM/zCuvmvTPUaPn8DH3OnDS
2S6JKEhnEK6ZqnvuudVeAPN8Z9qUocG2yVvaKaqiAFpMu/eej/Am1xhstnphHQjtmi9iALGqJv2G
Q8dyZ2IisvEWDSNwLUogeAiuUXgE2Nv3b51VAqy+TAxun09AySUGf57AEQ42yWE/gHfmiQwLrfhh
ASzOwEjZQGocR2zmmmpPuZqIPkuBH5Kr4RVtcNqyYqLLXEJnwL/gmaRy1EAGJTTEvEUBcSHoT/u5
pnxXJQAPYsG6jHgcWChTet76X1wUE/dzzqz8ubYuuSNw1JhBF0HfhTD4CDI+erPQXHzbYFp6yuTz
ZUuEZp9vv8jDtUIq2XvYxU9E7kSHUnnrpKc83Pj5/ycyn1GfG6+HfJ79xEsJ/sLtRN1TXKZ1LFUU
cumaHz+/Srgc/zgo5hDJkfaNsuHH138o4nuQi6hOl7WLsmKD2xGe658CBnkc7PWzF0axXCDo1s8h
tAqzHIiche3ZPhQW58le05eax3hcKmQdNL/6j9uNvtiGmpdR/YYkchm5y0V70TYE2KDXCJXb+FaE
zu23m5cYvmCfzbhPv9fjEZ+ALxsMHcKYyOTfPmOmdl/ajIWFpmpFwroJXgNpsQnxncRuHK4N+HSD
xbgYcj71SfF5bUYpZpFROn1snl3qv5/JIltWHW1zVlFRsxJvfea8JGF2FBiCcKKoiMhwATl/sO4C
kEpD4cYPBRFGL+ENiVm6oBHhpWvjgoH59FCdRwtKNNChX2onyBRDC1WESSZkFxRbIfIgHiwu04GG
jjPMb/jZpSsL6+ZvKvmGkWrNqTOs0miMCh//WvwAclfwoAVWbytE6wb08H9lSS+nr+uu7o/LUxFg
IxcgtiTeB/mUkkZT6adXNseQGomEPDUvWF5uNymlFdNicthWfjdw8XZ8UvWxwVGUlR6xjNJxQrJm
ZkUHR9StrXYHjauXGq0lyW/94bNz7jDS66umBTF8nvv/TYnmlsz5C+l4gkOTqzXPBut5rhZetTF0
kci1Q7RuB24aL0G5/SSzBHf4v+fnbprRs/dqXiKG0qG3fY6q3pwmRrrf3w3dkc08AsLkAfK5We7r
GEppVXoXa0NHHvG9FZpv8u/D50B48FnJUypdq04bWle6RfBoMn+cBtTuQ98k+jYciUcjMIH7tbs6
BJY1wiSvq+Cs74Tsct7hx8LRl1+uIT+18PJ1dAFf4d6+BmkmNnuTFeVufwyym+e/EGdIEVAnXsyW
bXRlciuYDT08SZSAzl+D6IzEGxX/UwhjM/fobjOFwM1FLMhO5omqNUA2U75cx9IUtWgoGDYUqxhT
fJ7m2hTkvHP5DrDShapZialAwHPp22xVQn69qWRbowAnljkbHQTwtmXZJmdSWOWXzP3lxKHgmuIJ
ZHWEof8e1SSvDx4vYL/G3S5U5EH9+M4RfXg0ojLHneKsSh5+b1C/7MZXWwPHqwHyKnJ5UMWsIheP
HBWPHNu6fzI1BG9LwHWeICaqRUqqtMut9chw4h+vjTCrNkUNpeR8yDdj6nOp658wpRxMvwIiT7FW
DMe4qVSIaRIUSIy3IicmKM7MIAdART0NboK3hgxQKw2BznCdYhYDrJFFhvbJb3xfTzEMK6m0z1WE
Tmv9ucdNtXSU7R+lN5xIE1Jff2SHFjc46U1BoGyTiNErMZG8T7NcNl/O3hqMkpHGxMjzXc0o5H1i
wJdS/lt1U8UailHY8w2zSRsW/0YHd+dFSSxJigcnfpOcg6GRB+FHMYl1BPt506roeWknnVcsdhtd
g0j0eHk+lAspYI+eOTvjmj2x0n4UrCJmrM+qD7ZG/VBTxUBXbSC2gxD1x0nmraQygoiDpirHq9t7
msrtcVd+e1fJgWrerzFM2wl1j8Nkgtr/1zmbgjKd15Ov+PJie9S9KiVNsVC3AW+F+o+roIpPbvTo
alGAjc5DbV2JoHKgCiR/z3bxJM7GGHBWiljl1rAfWPQniHjCMAlEQ/RHt1Qhamo4ZoznLDd84hF4
WeBmNHGZaBqVmyZhwrPWWnyBLfOzpMXZuS3h2QJJLEgZTA+AmKCs9CpkL5cy67BHEmNyg0ogLZ+Z
w3oxGlJciJqieDPFAjdbZolqKz+fI1ePOkYOvISts3PZ3YBMk4Y/ue4dD1oqYY37GDylwgt8BJQU
nrnRMD2qlrWAdJ5zfCEeXUbug1P4N4RpR9xBT1GslxDOLYDnTzvM5UM2VU4rhlvwM3wkpZhVD+kb
ZE7BFAXXtrPCe861AeJjvJ4YKx1v1b2weW4Bf4qLLxTQ60uxsROOWrvZ0MPuhJTOPz6derbcUL31
Rklbqg731urGgOPbaWu/FEwq1tvD817kY0S6sglefiYqnJmqSeVZUzPBiXdkNViCNNYd6hkwn+RX
LcEOz8XgSBhPsZ3JLkuTIM6Iaa2T/So/6CDBW6virifEDKNT32kNYWYfan8CwfQqWNzNK1LXWmTy
0v0ARA2imyKjcpjR5gFScv7of+ZIuTf2id8TheuNRnK4XzE415+4o+0jDBSFpytaEOmyDvMvIvMi
aqRo9ePEHz7SAGeSvFch90j+GfaoYWpK7wZQulebycaClhaCwIE8bbAnWSUkL5Un3+BsEqz0DbVx
14k7wYOS8UcMVpNK4ELnccvNq1iMuEjqs4xlNsq0ukgS+X4aurJ7w0YV+a4ns0fX26KMzxZyiVze
f2fpRNbWnWaT4oKBgJhw3y0po0GYigrkPmItFC/ypBSSR4paC4lzKDTQS9oSRzAeSxtfpCSwawFx
fBV5MgWcaI1f6AXehqboYKc8X6n7iHIYvVVxKuTc4/z0ycWfyywBvxCaiAoQv1Y22YQxjBKrErgf
FJzYmvnXhWSwmIsRSrLnK6JNtaipAASRSyRNT4BiH6VVmYV5hsfGFuklBmgOWX/mEnOSf0OT1PUQ
vBTNn2ZjpVOGs+1NRj6QaoZv2PoVjkj+LWC3Pu/qvxZkfqKndwQmYnQxitEBw3AQhCQlkwA1u4k3
vvg4PHYfdQCSHtfncBhc9VF2BnMCKxLMEBHbKe5IEqGRLV5GzrQfRuv0J1KizmC4W65DVFaePYG7
qPTYlkdb5DGvSBsUO/q87EnbNtus/yeMLalzGgD8C04WBAC9R2MZxt4k1/UM8ne/q8Zlgnm2M5Yg
eAsNJYgIdOTTdY9poMNy9d+CebQSctylHqniLuC1EzJEWoah4HDSdfZNGERNYQDXV+3dxzpIbgQg
gJst1aRNPWbgi/MmaFFgw6mmgztxyaJyQMqINQgWe4t3jjuCLjfyG40zajYaheMQ24dkX4ScJZ1W
SW9nE2ozXA0q7b0en/CQdFPZoZH+CT9/80P0jKQPfUqO7xjzwJLoBuzgF0eKPHrdstcbaaLojjuy
mn1RcVwbAgGtHjEuaVhZmIRjUyNCWCgZFKEddrTF0CzjIvw6GxHbcUlgk9A02hHXfjvTfVunqg0o
H0fHtwaSR6cKMpTX/sjg8lrDNh5SEyJdlsP0BF8Xo2UIu1p/nHzlwjA/9amcpYgXn/XL8kGUtTZ/
tq6gOGYUFNwTS7aMvXOwRIAD84vPIuvJm3kFmTZeUsRTrkDQ5Jr2CqYR6LwP0bpb5dNXY9N0RI/Z
O44b/stvKoTwMKFlqffVqK7U54oxkdg0a/diRVnXQUPfq6MhxdPYfm2leTAqXmqkoHUQTC/ieoOT
BM3W/67lgKz3k0yc+qPzCW4SOWzI6zoZDYsfRLUEouw5dbhnXCADrJ0sPANbe2LEIcSmyYUcF1Qx
YRBc/0/avquL7MrP87BY4Z6d7bJX0VuvoYXRC914IX49aVjcM9yhk2w94hvoFNZZHWN/NMQSUeYr
11+HMJIZMSiSFmszioIu6oxQgvaXAdTGHWwonO1dp2stERdpboKRcLUCnkGUz/5AjYUvlspFF0ib
vOaUTt+p9EP/oRZ6Q5draFHOzOKKzlRsHTHjE4y5FRKQjREA4+YG8Q+3fEhiA2z1ik+jMaheia5M
SgFJB+G78bkb0vMV7g+rUIKIvv/4k7oge2C/9tG+jK7GYGlPXo12AxJQDvwl1SCIUd8rW8LVIJnJ
GC/D111juvuy5PnLBGE7MpenS1WP5eNs3/vO+PaGRTCOXmOg16MK2Sc5dMRyn9s9AHQLQfbV5iqP
8o8VA3lGgcKdO0lRQk+NoNjvQfgGVOAUzUYhhYyr7omV49BDKU0WbrhXv9iFGOUd4kbONT1L2rYS
/dPGaAxv133wOw3XOGYfI/HSPnx98u+FRJ8/xypyvzB6MCX/q2bpskwj7JEkbSg7lkErlVOOFojK
wRlF/464bxGcBS0XdN+55fT7xVdYhKEd/Vmfd7X0q48Ozs35iR9LzG1ZCsQcnGxfF7pOIEv0mljg
b81PwguDgLVsETX8UILm9WUCd6nEBYm8zk5GiWxIqKwFE8N5CAtLMLRApbbdWIA82yQ8Oj+6TRev
LesKj7Ocyo+EaDB0cWieZISnMLlWFrBxQaNkTY+psD6RBnI6s44r1aC0Tmflih5vzRh0Wlwz5jtp
RDfRdvv67dktyKU9uhNCiVeYbXjYAJyq3DnG4eBqpUOCQqMdsXJBUGWojWZGvFvgm+r11yZ5JdG/
9OSzt1FnTFPSKqCJERNlAoNJ4XNb3ZJf3LbP3QtYct/xWhArhhBLnrOhofTnhTQw4er7k485n/i6
c2gh1u04RzfEXFUe85dajoqCji9LmZo/h2H1wHhdxQl0f13ej6hEuemGCIqCFwI/fEHNgc8Nvpd1
2qNEMg7tR28sGjPwngOFm7Xr2B3QICqqi/MeLgwoKFMSNzNYh5LCHohGtVbjY0pXOMrFCUXGc5yP
nqcWAMACmlkRVai4+l9/nNEjbz9C+1LvNQzvtUwwZpNxcwCENBli228Cc0k/3dwSGvCjLfILjPMk
wZEqJnPEAFEPsq1udFCEmkdy/hcJG9iFZDjmKs5Mnm31ZYJ5UyQi/+gIl3xc1LAmI1TyEbI5FNcV
nBtagpNJ3tsHW8jHTzM0UE7K7C+fDZV2TDfE3ohZxl9iSMFad9iziuS/1J0dtVfCpPbI9KAEw1Uy
FY5Zn8wqW2R8+B1maEdmT4WJG0t9BYXq4nFq/B49Hx4a8QZ9m9OSj93py4GoB5JA26OSQCwChOue
SkaQk3oIHAoqvG45UqibIxuYYChSHmjUYHNuEA3iOqCBN2WiBdauTM0fT5np2KWN9e2cQamLq8x7
rdifw4czlROEOPP/R7lXrIJEd/kWUGqJBVg3sB/QAqyt5Kt1ecD2WnV5Pgzx9amQv2rJ+E7xTgpe
XswbNHFp8QDl6A61X9G5AEfiI17X7qZ5TpFyITA4D6S1kgBY6GKpUsnG2DVwXzYY6RUvXql51uEy
fW3XsnamILoLcRT1ZxHWa60CEG3hCCR/IOr5wK2iESxeO3ndkgyIn32KTvZqyGZ67s1RFnoLMUUC
bysSiKDLhh9sorJVlMmuWoos7zSDWET9lUhyz4JBRvPtVFVABKFhud0g7OqYv2+0JKp78cbinUsU
39JBQvwg17NVy1e9IORxh2y702BRhXlXkD4kBl/KJNEEUuhM7MLf0t2ZJJDqhxjPOOPX8JyEw58c
K1+3M/qmQQ24t6uA4niEB/IlxdYn1P8FbPP4xzm0+LBAlD2LaNDHRJijQuiaZEN8RBHijZkdWYnv
PuRzwCO4zfUPVh8VFNwIrqHZf/nqyonyAfDJoEXtTx0VdRab/rP5r3bPT+1WV58DvC+0SazEEX4z
OBW8C/ScgaWrrJ2LT7/IkmwEoBsRTb+GOTwylqEbndjWVPf48YHNMKbNTkjpaks9/e+CsyyOsi0C
dLVBP4ZEmyaDO0k1P7iNBPAgIBgP94YUu9PMOmDx73BWDyvAatT/U9iLUgKxuXSOH0pt90nsbKki
fcJtz4Iz2FncaTELxjWtlnB+1hJV5AZ9451/n71pt0aBqFkH9LBEVxUK83g6rKYwluch+2B4nzbh
vX91eXNy+J09umlq5gZ/umT8xny8OlySm2CoaCDfUoSkyfRKEvA1JdIZH7dOA6WFeVf+0XNs3zDK
AJ3A9KIZuRMzubytbNcWNx9qbNlswVS+p65dNgJ9Oi/lQla2HE9oob7s1MLlLgyxWJreahsflz5t
jW4TUb34Q3Ma4hW2+H/PobJDph94qwPI32/uJOe/AdosLCeBmaKwK8y8GbECNNJPTVyaBnGj1/wL
RlXDjmPVNJTwaVfCPxifQkzW2FLjABEKF6BLiK439PqISexsSsaHtUR4HnhYIOMA5x8Qqid9rW5b
g++901JyF88SohdpgtHQNuOfWjVNDOSrGCxJirP0Nr4B+Cj3YH1JTMJ3AAEGisFhUamB4UcideWy
YLRh9Avx/AoLgCPC5yXCDQRRrHz/Pal5N04xvF7yUDNgoGFFw+fc0O4vV+JT/k/QLPiYrpsxR26L
RAQGUS+ttKXfprhyP8w86XS2q3oU1Kojx3Es1aU/RxWq92UHT7Qe+JikoX8NIhXwNV6vUdb4DiHQ
LwstT1MKeIx6WtHy4yMPNU4z3lSs+Monej8Gkj97Hgxzg8ydzuJE0bceGen1xpV/G2OSQpB6diAq
MdTuBfXb2vpCFXOTFk+BseXpZ6myiUZwEqmiav47549zvGeERwGgvf+uVg+nAns5t4AOLBwTPmVo
6rASO7M8lBKwjsISGwd092YA1x+bw6V4+DwrQbXbi6AthkrjkY0Lqw8fWZhioaIkWCf4LXSG9VfJ
FQ5x3Nlp+sF5V1+GkkPoYy6TR9g8FICtdPgZl8DzX9Y4ZpSt+SqMYQgwKnrasdk1RZyooo8qZeGq
Hbqi7c9SsDLN559Y3/Zopr8S1skzn3jyd2Oa4vvnSExyaVVVnhq19ukM5OhvrKE+rnAt0CXLZcRv
Zwg4ZtirwUmlHesApMR3L/zpW0ksmroJ3buhyFFtYTN3bzMmTi4c90e8nbMKpDpweC4N+pkh9RKc
JYzvFzSFSE7p6kodWFyMTXQxgLCuKi/FZZ34+HHk/iYrSdREOrN8Cx16EnwWO/+xxUeCe4m9enN9
V88ew/UbjGkT4dCVPUBgQrJpQ/qgHgk4oy5ISIPDWgbhJcJheRe1qX+k3btZ7dCeRueV1kQRd0bA
l4UOuiDM7zJOCBQnFCsxEvcqVrhUveTNigJu/w37sNtybO0XZZlFzn59fsvl5xaBL1s7MPSia0Ar
Y/AyZLhQYCMp/ruqK1UJXwjYNyM8JREQb4xeme6jpsjb5ROaesjB2YyCyb0EOrlztLGqMTwHcO4f
kuy/EQCwY5HwfXM5FbtNlvNe91amiDLfgPHOLEw4y0tUylt3M2nvi06WcbIPfrvx2kHwq/KwkDjr
iYjk+3DIhuL10Wl/vGK6XKe2tw6aQfNDeO9czBeLRwVT6s5PE0CSLejczxFjWp8f6SNlZU1gZzcs
AAKpeXBF/dCrz0VAlB/xtZuR5/+Bd2eNlqDu88eJMs+pYkVWVDIF8b9KHjAw6MKndOTV9VKAFIZF
HmevolT6zEyPLfzifzbyZ1+H6T806idNl6TuKwkHOrnCgLHJelkKYRl1rcgHXXoD7jl+j3jvl0bC
JdyfTWy12zQv50tIC9gn28s31PY5Ofp6DYJ8JjHL7VCeezVj9GTZrNCkykHUI9DAkyhm5n5Ior40
QcgDZcM/rDmfWME29ymYwMMcCC6/o9W8s/m7cm/9BJ3/aTP7qKq8FsRASYTDzW6gjAU1HxBvYiny
eBAId4iFvygaDIzKyNE0oylz5yfhvV8I/zOYDJo2TaYfi9Aof9Unu+q3pHHLZt+1rRses9pJfULU
GNZ38R9SjlkZ9kSfulfgumujFN7RvEMxMzGFXCq/AR25L5hvrSVpIJE8dLwg5kvvaSKYxOsLDZ0A
OHs5P4c5vLK28fQnlJjk6KSLczJqHt5Wer9cYTqBcZz2TCZyDv/bhyP1NKf0UDX0QDLy2l7oWGVq
zNdZb+GsKu0f2Bo+X0E4HFR2jp0KIzzk1HP1ihFS9uWI6VzkCvs1Bomi4BtE1y5RfkOzCZEgwary
JItcO0v+SHQQka2VtzS6tHmi92ndJp3qybde5oRqCJf9pSw4p6efbyo0J8mmS/9q9PIfTSbnjUgl
XiH8Ggjp2Fc0g87sAMQgaS+5rCuznW/nRefd7LwZXL9n+KwOCwlu7CNaiyOfLNkiRoOBTue4G3K6
Gti4TxqmWWpSc/Y9ZpmhnC5gckvxY8rqENKMhF3qza33rOH0isAMiaOfEuLvKrM/f4uwssOPDIck
PD8k8YwQ/Yhh9Zk7nkrihkkt0rRpafbAXJXYwTEiwkmWunzUJgUUT4fSyec0hTUK/w17HPgwpu5Y
pp9lw2XcLuuyu8tmlnHj+1nsawZ2SQ/qHE4dD7yYVbiS16aMQwSNRWn+t6S8+p6uNB73J5Vc00Zl
sQnPjGIZ+mKMgaKpwj2ohWDGj/gZfvk1KoS129h+XwWkVZA1DS9vQhS7DGxjeJZ4LY1BaDU0w74F
gtOxhdHyLUYPGdFiTLOxvgNh6YFASiM8cszitB5fiU2tiqzTZ/jjZN8bX0maJfYbm9KQoidVcIG2
tILdBdk8rJsh+v8DJClumsOerrLA44dORWAO1VXrTVWE9p1yT8zDgHOf+hlaURb2GQzeQouqu4wx
2KRXT+XgVQhS4uFYQkp+Bux+Hj2gp2T7B4ad/s3Me5sRUtm0JKLoGqoxKPTZJajljilE3PiwherX
ydg0cCmr1cw/tP92wW16VysCuTWPpBJ1+aFML3+9rLLuVDD2w5MBYXK+uBAq88P8LFz8pY76tT+I
9z8Z/Xn7suT1nPDIfTntEyBeJfrhyKD0mPmP74CNkhiqYDkkFjNCRKQh8nkK2nP0/L3+30FyAfM/
h3JUTB4jbqXGAXv4s99LAhlT9dLLnf0yFXkhqPPe5/ucWfLNttHY7VPdKTWAfUmCz4dX1B8DAluI
Lq+gMItJgF8zvP0n+zpJ4iYMzlFMwoRFqu7efIHFIkWHF7DNHv0HxGJkG2wKA+2jQWm4vbj2H+wL
f2241cpcnttSQXGflpqkUnQV0o2iNcrvRwpZmNQ7iqsPebhasbybZwjdRnR/DowsiRHXb6lLbgPu
ZZM9G9AwGk8un1s0ohJKsajMYesafiBn8sAnCwbJNJTtMj0p2t4EC61GFfUh/IXCKDuIU7Ae8Oz7
SW8fauyBkzPfoRlnwYHaZ2IJ/2YQBe2ghN+CpXvewesLLHrpobV1aO4+jcBIZAHVZo1c24cFANj6
k+yjVhq1rxGQZDYHAwAS4mP6lHZ3wTlS7T251r2zH+aAVBxzb2pX+Fnfs7Cc9yrVmEcMlSeTgYl2
BX3dG6CUXnTiOQGfyhPRJAPmg+DmbPxkVk2wcWBKcg7buHDui37lkgOispoQ2NWOYLQM71+Olvjb
Xj4MYCkdqRnEscjNvJuu+l6nx8cQgBZh0bJD/SpGUf/qH2DCfXrJAjFLRTK/U9tsYqTDFSc6U+4I
wkaXqU0HKQmm9jpuo9bDWTyrqsoixmg4nJxJK0R34OLVZF1aLEolnnWJffGM1yf00dZqFIAjg5C7
kfDy13LNfs53t9ivni4oZg4n2s3tlH8W/q6vU5YMd/txzubGvYDDmdqlyx2XdGCQnKQ0W0RD5d9S
68BWEX7AzERJo10i1rw7csy5rrGFOtC+bQEhagFPTqFtojzKSnpPVvlgKv81oqdsrDNtjBp1/+zx
07Af/pRzIPkIXZI2C2W3CfYnhBABSTj6k35Fv/dpjflhYukAl6niBgZhIzBejERIbX4DkPADnfQ2
36t2rHHq8FP/Z0sWgAs4YP388ljtqKqv2GzjLy0MSY6aVVlnOk45o50fGRuv9pPLri/wHWGH7x0W
LB20scub2/d5EfcRPXFxBX2wj02+77ZfjoznzvFzjO+1tu+WbHyVQcwvw1WMHpiVJeOPBVpPpDKh
fH6DnK2HF6QKSbyZAWJOQoPNkxtjVjcUX0NdHoxhCrrMOzwOJY4HyvRSTmieLFIAMjTO1xKBeZbD
jAHrGqHjKrUsI/gw6qYYx0uUTsqjrmVICvyOgWAwf/HdzgpGU1gEgWaWGO539VxkmvZUzsVn2Kyf
Lh1SQpBjKD1zHHg1lKj477rWsjEOkWL+SM+GmTikczN9EyzlHIRz+R8Vat9piWcYWC5cTqqOSbei
dYcYa5UQIccFYGRgRFgYHHF34fsYBxGX3tbKam4xpZhvHZoLTUtXxRFVArYXG5ZPY94BfpWZGbxi
66OosmtLcdgBwrgspEhf3cCqeaMxfiz0j91z895nCDhqjflexulM+I846N8uS3vfQPWgIaIdulZu
9X9G53gHTJ3hPXSgY17iS64iOVR2ox/o4f0AeW1OgwwaWcu9+O3VBqXsVlfFYVSX9H53n6KYUWy5
AG1skkzTytjgfYsxqs8Fm1MsPL24n30RbLVxLSusdASSf64jO/XmNfR7uRlJtPdymqg7JvgdPN7m
Px5nZN/EJYSHkmYNepgHssNL91YCLSrWeO8zyDmnXiTusIoip818fZ19h1QUzL/fhuHJ3KI8kdbI
/hw8kuNi0WNGrjlK0pKvz4OyQ4iAGTqE+lDSeOosOZJJRQ0CGHg3JA/PwQpLPQ2CyiJEomEU0Srs
U6+hYjnUaHWV/2EbHrVSGiVk79yB+8ghU2EBytpQn2xmrrMH6Lm7NhywdbWtPcxTBy473sG7BD32
VkR0au8URMKkjUc9jIfZbxjoqUR0ben9zMd/cknzWuwb87SQJ4UVe1rqQ39DOgHrYOdqM0u8QGPl
Y5xnwF4QDBLr4/k4BPIlIG867YCjvntFrZ5VECXMdbeRKZDFfM8RoWuBUhtAzqu57zJihakc9vrp
sKtdGKbviiMVQpczBiNQH9jU6Z7w0GuZoUPDF3wosLiu4gDyrLV6eUbDymfa0xoLzno4vRzFq9nB
vwjOybvWMDJNEbFj/+uqArcWfvMKnQEaFRhdjx/CCCYUk6SvZ0nKX+/ao0ljUaMRoFiQwsvdfg6T
m7eJDrBfcHVvawjtmuXSsLdYhlzXKy9sq3S23LBzln+LUfmMVsroLbk3KzEBX1lQiQogvHuqiDy7
BI/7gymrLlpop1y+bTSZPVlB6L14MMkBnngd0MRAy9wOXAGdaCsf4SD4xhr9/J0WPwpnera8z+wB
V7ICKfyufyEZ63wA2xKo7wR793dNAx5XQXvYjFspkr2/z2Bx0jYfykpTeozxjn51G2KgicPAi6v8
FK8ASPGOzLHlWGktDeKhe8dmUDFwVpVgzMgvfxT8ctT4B44FcS7ORjIg7AhhLe/DwZ8C3I5k3UYH
4OpQajsk/ey86jsJ9mqguWZF2jXPVyYUnwJmrtbROOxUKyohiUgDGZqarzf1y8nwHZPySafyHkNy
rk3SQg1rDNyIwyAspTDgD8B02mAlUPaP2SBAU4MleP9IuMfJ+h/Yh5wdb36ckTI9kGzEA+812trE
yNArVAdZJtxNHXbJ3ph+1eZSBBbZnXsWohSiQR/krvItlr6jWiy7/HopQpnTTsDcdVOW0vY1AUrH
NP+6auB6g/lc3eTkYF3DCy+efcfv97dZsEFhaszGTlvn5YRh8S02Imkdqf9j1uVuXdFQuq157FS0
buXf74AJoBErjKz2JxXCvAc2+k4kWzSJdT0mEhg5hJ+iq01kOZ34CVveQ5PFS0WC+c97wfqy77OL
xDSJxf06CJE9pENB1nHPo40IPEvdfZZjV03ABS7KK2+My0LRSIW/jXRnTKv1Vt93978pSOTk9ZuN
u08JMQbQk4TaYZXYM8BNjBPQ5JHfGdhovTM6sEDe1FrF1p1l2mtmY4+Q85mFpnuxaGOdFUOFVbrm
WsN/su5Ug7Fj5wxOhggAeq5ULo7nFr+QXtG4rRQNyZ90f5mOVpcn+hGrXxa6wKrdQorla49OhRiY
WBU4mQkdwdVqhEODDaeCAtB1i0RwazJdpYh44pq2GDtB+t5dY9i7c11I7+unyri7q6olpvfrRbFt
4UbjP9pxJlk2TeoMjdScutJVomRNO3HLTxxvHfgPdYIYsLiC2N4fjD7VeifjPhHC9oxEwITzkGhb
e5tFBUjVc6lmpQjBccY7d9yLkVbDRqu3sNknmjcpFEZl8auxuoiTp8sYqpHcdPy3L+p0amuoDJtx
M8saae9erIGZws4RajTUpwrYLByaibkpHp+XMKwxg+2+xYIUVWix/iM+5Vwxr5MOxsEMu5P1jj6r
f8b8/T9ckhebg+Fm+naY8p2p2g3/v8LC4HOxr6NbU6ppDO9tOr/MUvBODA5yUGMqVqKR4O94JH1m
XcCEY1q3NqemVWre5PjdP7n3Q1zzHtNTLLbYMNIknXOU4PzkFNQ7T3TSEZrmq97HhZ7sabq6JD2D
PG8w3ikm2qK8Wei8k1+INDZwCyVcJzvm6HuKXbuUSLNEIwj9jaV7OKQWpvFkg557N4p2elwz+DEA
R8jFp+SknYPlso1Tdh15+qI+k/UJJtHrJPRVUc8J8G7czYwESihEoqWaLf1ZjxpQSNWOrkHfSRd4
gjr6IQwVTNRDHFToQOany8U74OswYwEui6SjgsH2PKRqOsQvs3IM9Cod67fDJxQV6ZJBms2z8EMY
Wyk4y2tUYwnq4pQjSD+dvZhh53RwH8Zc1NEFbKD4lI0IEwJmu1XNfcmdlC8bscrQulI9wGSi/ylE
iJbUjfMtnFfKIX2xOLHj4onOii+044uXvUbFM6nniIhq3MSdlDC8rStxjo1h6KwhsyWqWAR3azjU
IYJewAGtInE4/mOTwT7efcFgvAna2gCHWKhzgjFpQbRqznAgXPErgnvuamFCk9IPyrirSvXhu0kP
79bU45ry+0psnczV3FR4VrFG01Enk3sFiP567dJ5gjoDzEb5Lz2d+yGXlbSHdBlY55T6VjOttVfm
JAOaWDn2TCmW8zlLVhRGK7N/1FLcxbZl9Gb5WRX5BnigEKx8lQmxBVjYJgL1KfCA0vsoH2ZvNFkQ
BtVVOB8fKIU1BjlYOEEUdxSqspFsYTKpJ0D25QtwQe5dC8LIWWFuRSWzsNHBic8FldYEh++p4FID
8ir1kscg06rHSqSTNnsEOaKGxD7y8gvU2ijISJizgyPJ9Uvb9TfRYA5TbDb1dowzqItHeJCydVoF
ysCd130jKkuUZ8JNB2i96HtYYeZNtxLYg5BHOCYhPnL1UtPqA8kCwG+h2KKJWoWS2zRlXZrPzTp7
vaZxfvi8+Z7mfQtBHBdZtKz9F79CBmuJiYPBxwH11g1S0t1yNAGQuXe9V1RThxYXRxlZXJ+cgNbV
e2/L0nVrgfwc0rnMqDE3ed9ii73D7aKEygTdqQqdWU6Hid3bNei+ThuEzS6fWjg3n4TkSANxbelJ
+zvXxpu+77GKi9e1ijEr94dt4yGB/qS5SX8pWWNGtk+97EUwpzIfq4LrK9XVeW09MFMZSc2crxPI
gm6qzFUQRNfYBRExIQOL+qrojgmLu9m1L1LisElytfKZg7SrQRfdEaAqCcL3WTwr1cuAH5EjuPzS
FJFvxpE3Y7rZa3Wj6/kDQAHc5CMcRL8z+fOeY24iZQyJ2oetMk04dcH8ghXfYuRMFgrrlLsdKA7a
4hDjfEtUSe0OQ6etoDkASLI6EJ9YyaUjPQXN6xU0pBHCvL2t5aZCHCF5rdpXTDR5ay+TyRXBnY2L
wmmLt+1VTS1USXfUwYZgRuDxaR87FlLYrqdPkd9sq3AXIADNjO4y2WeviQChvM278umz0f0ngeV1
XcYsytU7mIexecXTLSgtzwt3iuEFu2zB8WrrubxwRD6XZvP7AH+MRw1NSvRjId48DY2GImSCEIgV
KRDflceCQGFG1TpK1Y8zdoYkIQ8Zy4SyZJ2H5/AhgQ1pAKdS0e3oRczEEOUFDTe8r3C0WfCzeXzV
CyzshPzLZmPW0Mhl7XbGo/jfUOXe51ljnxBfiPart3/dbNgX/atVIYQNNMOB9G4MP448mSzARGsq
LdCsna8FsyFhba/5t8UocBrD8hSjUeFZ/ofQVa4MOmXNQ24COCMXuenR6muNDEkwKhHXi59MzIOW
P1Cz/urO9LVOCd2ntFDzpNTvx7xASXvRg5NQBiIWIQlaYGTq3ZCVfNlYD68RnjP7Q1oxuCTKgRxl
KDWALZqzY3u1r9M3oUD1y1Qi5BjAzWIZQd1Zk7Bk6rYxUHYqMIcIqNWrGqwE5nSUv6ZpRYMhSxd4
9czHtwsin6UtMH2IiQfpQbS8myLMR4D4BQbxWk8uEC6q4pWfJkhS/XFqIjEuXfVXxI0uJmzkthNr
uM+jjxyRq+q6WBwKswVVZm+86WgEioS23K0ZgNdcddOI6nnJtkYxuu2i71vjMwkXro299oS7ptMR
OEONt5l1XtYGZVlNt7IGLPDEwWZ+vv0mEjMQzlzbOOYNNNZ+hpSjwIg8E1OcppYtBGwzVqh8iXw7
yyF4ivuLfk0UhknknOwzf5+yB7Ob9jEPg7W1/rT6isQ78odheNlhcWQDIaiAklkqmiYT9rM+UfHD
XKwyI3H4roKVrHueBZNSyd78wPZCRVbp/iXH6RVXPiWx2YtgXhwel/6sUzihfsJu3ZjpIU7/6wT2
KnJNqfYzLi9DmlTB3WaZiNgPOwj3Sx2m4Sm2HmM82IOFpGmwHkoPwMbcm5EM0WCl32yUaZx0+kHG
j4pELK1adLVk5kT+rGjl6Tyoh+XDtysdlfl32xuzbZKNqDxuPb/EdvnmNvau5XusWfp7MmesLke8
HjIkmEf9nkshsNF3jN6PnyYdzFYAnvl3F0/OlWH3nR9RUAQCtMJuPXKYkzqSRBDC65frplzWeNzQ
aP/VJy2fN6QEiutilIZS7Acl9o4uj4NCV2O3VTVrOsymQpVtmfCRgF+mHQaeYxpNdctLGG5YEOml
/fYhB6Gx3FJCrKlFGY2giauHOdIwppNLYtkehYluGikpMKr0KJfwP6IxKw2/ifB/L5qDbmiCywNK
7Uo1fyym/xaB3Bz1Fi/f9RoYs/DnpPpJUtYuJj9uiuJwbPnaO/nl+8s5KfHEOFQqy2vdGsDB6VYv
uq8LAx8h3q79OMmUOMDC0s5aNQ1vUhxriXDOEjO2iOk9pXqFNXI7s8HzhkWUTMk08kw6CK01B6uc
VFqRXfXqGPtIzSjpBqsI/0FotDAyYCdLmz4uOrwtAKhuIs6WKUtXA7yBC2XmqLB0SGWKi7+lIkZA
UYjDLVGAFPApUGMD0zdqLNWWmUJ7YiD12TXQxDBglNSdP5uYw5qz0DDI1KzvFjTG+0b/BgMcx1yv
UyEQK7PtD+x1yR40ZHAQK8s/vmjqB9EPjFHK8XrdODGtOrsLGYmJPKK0BPZX17tCwd4Bewh1jOuf
OqMGcrI9h0h7m8m4KhHzzOfEfhDletVomeUByUvKfe94nmqcup16OjNjkI2l+YP4zALX7ElAYlzN
nJn+aB9+vXPZSf8znCWjZeiI4btBunld/sEUxagtzLPa2pooQEAcyjiXS/ow9woF+/uh8NDCQCPC
bdQ8xZrEhnWl8SuoDzXK4pZ1eJfbbCHiKWQ9TIrF7h8TiaTpdjd4EN4VF+vT5llrraBYTNini/dp
4sXTaNw/XjW1E9vEgg4kqtQeaHAxhHB/lgdnBZTnGuhzIS3UCsntV6eSnr9RZZn2X2cdvyQvMEBN
0hVTW8F80Q/t/jMdow4oPT9CLDto9Abjp0xagzolMdJTL5azxihqbOy090mYvRC108BMXcMHAkIs
TW0eoU859uQr0qd5ARA7QtiwP+zNUp3AB1EmCG4pw/aJ0dJoAO64XVrXOGTxq2E1q0CLnTvEsu37
FS7lNzS3pzBnk5cLStFZgOFx6/IcOylMFv76GvaL0mNgjuwgQulAgiYdoFIo6r8ysFPiLi0WhQVu
G53hdg0/MEjMbPNo5C4DaD+IGOvWKS4bFtiKcDFuBvFYMWJRChzUwXzUfaHnrG9ezEF9iOgZOoxZ
jVDgyr17TxVyQOBK+Bmd5dnJ2r7loHorcyWmJJTqsmsxEks5rYW9xE/baDmw8yYMztrY+euisfLo
BUwr/ye91j6uG4tQYdnUT9grDUw0eYmX10WjBfPR9/oCNV5CiiTPuITTYQaI+C5oQRrlgD2Dm7tZ
tOXAFhHRLNpp4vcznIVdbYyN5Xj4gI/s6Mb2qe0A/+lXzK57X0SWfCEsdXfWaaDHZoDmRoPm9/Fq
rKejaF0MRHUfl7/8Rs0b3GEbQ9YVeUl29YS06EnZrSxJE0JS/Trf6rlrj1ePA+ruB8R0kN4KXGIa
qi56iTlFlGZvGhc3PVjaqIMb/Q4bG8kqSF6IEEMyJhyOweEvhWOk8jtAmxaqwqnnzrOdTNps8o2t
yvyxrNK+UeIBfPgrclnKyHLqh7SRquW2LhSH5lvTQXiUxMy7rwAyHp1Jb9zXtQlZ2+mlw/AQFLF1
kCWAbCiOiRtxv/xwv/sZZyJSuRrDz8keJcgNOrErcv+P6IiKj6QV/s2yu5b/fzwcuVfYopnMH5pA
fvsgyJZTB8JXAw4O2d453uwdFebejKbzvLYwMpmVVogC5yLPhqCkTx0jgOY6xoJmZ6CWNOTSvA0o
I2qOhD0ul7Iygt5PTq9xJGUUhHGhI82nE23tTRdDdKYHv2Ei1Kuv9/+6fcC+OXrLrFNFmX+5GBi5
tOHyNRhHHDp4uIjII8QE4E5uCC3XVqzB6eyUAyo5FWZM84qkiz4jt9IFpxonJfXxaNhFvFbxZFBr
BRNL72R6CNeb8y1IshySsF17AS/o+NNhK6kIymfW5yerz4zuFOAplCsdwvLLQs/bQNoxqOo4jveB
1kncmKwA1JdCi4g7yCn+hoEOG19E3qYyM+RO1N9uUpP5ay9XHyurwi+JwOyHK05z+1HudJa6YpL8
uZdvwdvfQ/zC46kKexUjYMVbDCaAHO4omcJjSaizYkV7zyPqHdp4HuANPMOEgqjUGJT+NN8YiT2/
klTTOaiH0PXpsl3BXfiYN5kK6bKajf7L5sD62JimSFhVdXZFlYDb/nSLXtttPrq6NoKkK6iQqi4g
rhgF8yDzxz0Kzi9SMf2Bb89Rlsf4gjp2wacToKpZRk9ss2i3WSNLUZoXytpwTP5ZTylo0mKKdaLA
0m4u2I1C8yOqrk771xi9I0eSQj5csJdI/8GRltst8aQNp24WEP3nljZvNAt3OT3R9I5KKSvclmJ3
APKtYWyBPt0Qe94b9bmh6zLPBJQIc/5rSjt36KpPWnFtO/Fdx+/Iw0IeKzaX98JSHj/ETKkLeh8Q
8X3p5X87JXXJPDahdf4CXR5dj+CthAdzFZbzQLEAFVpTBNJCQLB31jvLoKjfxzO/3blkcagQDFA9
H4fViKgKGD00t9M4EMauDPUfWL/lQohEp8y+/BnijOi85xL68d/udh08pfwrc2rwVmx7peBAi/nR
bggO9FKXltNPuZ9A9ovWFOWyEp4TeQYOqRFX7Utxco6nTbCbw8la/WlTvEQg6liFCni1CxB1Kyp/
PyoRRAyuAf9nywJyKKuZqHXX7TTMDj/HGR1ZM4/73sfj7T6TVzeOqwH1eqJx/bbtQjaAKCrMGLZa
gHqfNnNbQsBTLfs9JXgNPzb6hEZBkeGjZ5R0NIXcLWllPMRguubx4uI11RCkqmCFmpfhQ4/w0XYV
uRwVF3cZ9dW8qHVG7W7qv/9QXbyKrdjJ65JBhRveh6ZYytXsdF3CCeNrrIjto5oPn+qkpQ9yOAl3
nhFy5WCnuT0Ptx1lY9jCgs9otGQAX7gPZs4/4KYWMMctnmVqFbPnZWNwxPA9Yl42GggZVmPlpkep
7YSM2gePG2r8e0+5U0xZd5iSkTnJpSTOiXJEI8vnqaCY4nHAbLkIffzB9rhIwXfmhFwNnKGawLZj
21sYEio0WhGYzn7FfP0FHc8xSQ9+H2C253oSb9WoY4XzV1Bfjj2zq+PhcOPH4hB+br1WRALA7jM0
xPfUJDhJkTdrLxtV3onPw/WMGx9eLJ6xdxudHWKiu+bA0YyhWJjWieHHe818mOFSAXMYPgL7ySAO
UZL0+6ruAI9ObneN3rxdrJfbcGZvPER5w2n+zoTyG/AoR98iFpRfu57HFUgHYlWA46VeBfgET2er
gXgNizs4rsspd6Q0zgS8ClaKW2UMzHBzWdWLk9yfQLiJ02wCs9ukDBlPFMLVniw251olOKsNpTmt
ldMCtifdrqR9luOmsu8dgDweBeRbcWRXjdiH1swsc/axAdSaq3awNaCMgIcEtRIB4iJgsI03q4L9
xRxTySGkbQjyFJ+b2MZOgssFo0LbuXbOW2t0bYM5SoKWq5kURmYwgKriP/Xz6Uat4lkv8WBb6aKG
E1fHs9CFYcfNyhNY10GobPbv296iQgCjpt3SSDo9TLIcekAFJsT4hxdiwvXjsH5EM53X4N6bkDyP
RAVvJUY2nVGaq9cg87DbECCftzbNpdC6X3MtUXxYllM3V0MPmhlUCmeImRKwQLiANjx1szPwf8UE
sZ6RHBnfJ8d2KaPdvWH/EQUS4xBGnylZaw4+/XLPalZTnWFFrzG67RPj1CpLnnuIvTR3T20I4Nks
E8kVjCG+3qe7gio2N2Amx03iLKfMI8rD1brbjZjvhDPjZMfGox+xhAoK5clKG0G1w6HIaMVM7CdJ
Uv0k3tn6eInLd/mwSAvGcCehQj4qtL8LNNl3PC0GSEsQqaTC0GVKrK8Tf0IjVKW9aWaffrGctG4O
lT7SlylSwmMUVaqf1asyrkM00FjC6SljIh30BckhzvWqVCcpU1CY0Jm/w10uGBOLoPuVR4IVPRb/
XIw2v9qryJzQ1AkVCoMh/bxLNsHnHOI5PVfJIgnmtTqoxkfsmc5B+1FmKaeRH2cdwjlBsBWJVolj
hvYESH1ZbAZFp2pgkxcoSZvKigag5PRC0cIlgSAohiMjENnIjwbw+BOy9cxn7hezozqpBGIINu4+
jk/zRDqvFBBB1HXsczKKV1OJJMadQlxYy9oVSz1LgUFiRE8Yf+hI3UsqGroskmYj74MscHXmcuIo
Vlj412e6lOngFt+Ggl+ai+yHQyGJ5IHfjCqN/LbZCXHRH0jH45yfdvzUvow1sRvWmAs991SwWI6K
hmYzBexWrerAfa0TWDRAQrfHKaPoyOfGJGB8WPrkAwp0ZH/XAdZ4UUTM/2RhEQIkP63yfBF7Hg2t
mlfABrgW1baElwvNneAxs1SUYPcI/0H/mlb37/5qWJTbpxBVmWhyzlXcF5Hn8rIDIK4aSxAEebK+
5UlWnT8q7XqSfKfcSlC31G1nkjdGypphoYNUOko04xBDkCgTEaAFXU9hOnNQq6Vo9nG0AfDFt9Rh
d+BRbFbZB8bXv7Re4YC6CLmrasYo45KfqqK2M4ct0s2RBFY4BaanLU/KcC0yKocp00SRgedVLIvD
otqWiEOylxt6PX/m31t130FE/z9Ikps4RdV0g4NXxlpy3H+Ty4sJySH9VjTPQXlDzH6JdY6Ryel/
IDLhcQDt97u5TkiccPPyiaZrRGhI5eZxrIdyaLroXHLSh/hLu65YTgv3k15ZIcMdWiGjujiyEXhy
27jMTWraiFORiNapc8NGppEN/29hsdaWRDZ3IVPbtkHLBTjifz5ech3yKsxtwBr6Bg9KQKWFNDFe
kxl3OlCjAaAJ3gG8lrDRoEjwiV7fFXljPgozwN87j5rZ5URbaXHdR8FjVRBAWXVvLO6JNRnCVJ8h
y9642bWfV0o+ZC8p7RcoOzj/3r/WKp1C2jAEWKLo8kqbVzHH7zx3nXxbPLopXLURgIn5GP/sLlWb
WAtRw4dH2UmLYNTqRKEbG9b+CnL0MdmKrSyQMqanXWYjs9ZyaYW1OwwXEsO+8g7/5ehFjZYMiOf5
U+rYdJXu7G0Wxf/nJKyE0N1qDjsAG5UFUFJE1ix26BmEzDJJj52P0Rqv4kLIVjghlgpz1loOUZaJ
6YAD9POva7eN5sd03KTMgXJN0BXZYGi5L4GeYLEEWqhiIVMgFHuPvOYdBnPxAYnu94seF844AKpX
+ash+wBpt1uzpCkUgB/FZMdTouhlusU3Iaw3FCbeWoceWMecBvB4fFs5IZ+/l31gkbqUTfhgeZhX
Ecm6CLR5Y0zWAquWhHDtmN4sW38PejKtAcI8/lzyuAwRpCFBubfu0m/PBPp0a57NurdI4/LgUnuj
CITBemEgf5CcoZSWyKMB9ty6hu6EYHxiak5iWLTYvF1z8otcawAS+VZLMCy6A4i0ihK68W2pIrYS
BUJyzTxnvmAblYgO8LwPONFDkDLLsdtWtGMISNy1fUeu317pi8y4gyQWnllN/N0gxSeWcXHlihG4
CjrbdM7U4bGhvlryUvd/tXwM1yklh1bFh8fHf5fQYZjYvAafNfwFArt909ZC8DyPgiyqxwB6rrmf
gJ0AodE/sVSqdS6JIsNc0+HfukJ689IL+ZK//GsFt+QglN/bKCphqTLZ6ngLzN3ZK3mCs/tsKlDV
OeLIIFhkEBdexRa5oZjoLlgUFICMXK8C2yTcAbYG5hwQz5NhucAHrodyRj/UZnRoo61nQUiV0otO
zyBp1eDf7bET455zYUJQ0c62Azom/8cUm2bf3ecpeg8yyj4YslDjvQSpDAYgw0wToc0YAa9Vsocb
JeMEfltyDxt7CJuZ/kiSYIjb4fSWVgt90HEw8BcV2/PV02S3YzTeRHlJBo7i5B6O2hQnXpablGbD
9w/hWr+09xtsU2mpF6HK26bdqQgpQgVK+K8HXcKcIFBVwOXZqgVSFQ49a+XNTfH8weWONcV/GS11
J/FfcM9U1eINWyFZEzExmmAH4fr1YRQYa4UTfS+ju62nEqxTM4wRgdK8N9mutGUWoB5tKDa+jHV8
WcuO/w90TVzDM3uyuwl8MUFmOxb3iLKP+VvL2q+t8bGMhQXl91Va1v2bs3aDmodYyfcQ8sa1+lKo
iEr4Vqpz8Lfh7EcEcGt/BOAar0qC9YiqYxgvqssTv98Ip8QYryNVddT8PRZ8l+JHFvnZARC0EUrR
AA1tDyOM+HaNOX5COglBt2qr1dUhBvKmPrKcdMLeDaGZLV1l+Jdz+RLM7VeKuwbKF8tfWGukFDax
9RXQUIFvRMt+d3DwGYsyGcyG1IHKyGjwkYOXefQki2ilQir+EagnkYxD0ULXJiGc2FxdMq/yKnb6
jFF0KLvGL+zZFsDXsZRymtr0latbNH2J9GSV9AA3T/mBCEk4pm1gzDkHXpqsxbe1Bl3J20MxiRgb
C77MOc/slrO7Tw9VvYj4gdAMpeb/zzpbBwJvqfVc8a5q5FP8yqR2rlGxaC8+7WwVyoUurm4eQhnw
ad/4v3NsEoW4Ay0RNhoaeA22ygdkz4/qGOQeECM//grk4YmFyW2C93E2SrwpznW+3tAx12rTKrAW
2aOfs0BZEfg3gM+aQKSgce21mbEqijwQ9iJ5a/k4XYvITvEfQwBNVZzv2t2Kttu77tKG+qqBIzOB
m8YMduL5VqXTMyTMS/G6e3eZ7owidlLwVGS984Qo8NpxI8WhOxYS+mRIQZmk1/y16QdplJJZQeXU
QzB/hf3Gw2IeungSuaWkUVqtWBGTmo2oTdoaL1uicf3Q7l8WyTtdsRhTbcFLdyGdhn5/153pzSNF
HrVGJS4fmz0Bf6VFfWQfEjFnB1Zus+9VlLE9vJlZYwSfOxxeRrccJfrvw0/SMjcTLBcMIPBFWQpW
ts+nrSQVt7CeW3lx7KozldSe+bSMYSvqICDOBv++SPopKjI7cyrHjOoK84uOAM7fGRwucbscTdqf
Ke5kDatO+tFhdoQhhMN0w3ZT3NkDvfdP79qQ1/AnoOwqooUCmuRulQ8003fVofS4TXyCSLlu8+6E
08YNScFF/3/yOYUr9FGw71RSqWQhh/ibtePObmS1L0ugDyL4tijaRKN7z6x8h4+yO75CZTPgEzhS
XVTZDm2BnxkoAb37+SwP5zImavK1j/GlmUSCQvuFIxvMWCKWOoYBypbAIE0HVTclxGYk83jwHRmJ
MnVYPuhEJUZuc7aFoFTWCWH1HMC54rx77Rk9WJyUIW+b87RqjMdEeIDXpI3gUiPNfieG4fyidpf/
W3hV5Aru6iNV4itknU7OGP76u4JieH5sYMFK45nGiSH9us82AEmpBDeuHs3YNh8MIOZOB97reTlo
o2Drdc1LWv+b8R3Mw/mg8Q7JJFjIwTxe+C0N1f77YW1RHAdJIwMbneR1UasoVQEwa6QUNMZGBZIr
kopUBitJiefGW0hWITBNecFy5uyIXhr4HJF3Vggso/HkA1VC6NeJJfe7sopz7rgwjhAH8dL4NAuH
18WI7IaMTBScr0gRpa0QRMPIvQTSMdvy/xplA8b1jqHCs2T3rSU5+XLkacehFva/iKcyFrwPKQk+
+fJCmOlbqwgG3w5vgaSyoxB1ZxWeQdWWwWluV8Msh4O2yGZy1WtV3IrY4aLOgTifc+SO4pMnHjR5
ekwxn4mShmDiB7U5BATfVcT4DFSlJ8F/+t8dqMSVe6iLdmthOQz5oclsEnwVf9oO3Dh6lfbpe0l5
UmnMuU1CUqqZnlRhq43B61g1R+GgXrXp9Av+nB9nl1Qaq7q4b1N0F0xLWoEWvAUcRv3Br6mXaQZz
nWW7Lxc7knXnXk+ufx1A7z2y6nV19wWDf2zsGu8kkYD235QHp/3bQS90SNYTCl8xAGIu/AV3BxYx
OlrXzGE4ddfMgh77TbDOLrwvgawituc3uKA8r3WHwquUxVame9YibCKmEOHXjdKZgc54zBrCO7IS
LeyoQwPJdQOFBud+ZI70M82+vWEGdQ3/fnOGsvvHSPh5gk6VnwztJ6vb4fUv0rwBGF7/StwoBaq0
AU3wR6qMC/8m5JWtlZYxixrWWXEEZQTMrJ9xkgx6NLcL/zvomwv9SacEgIC3r6HKjzdtDNCZiTwS
PLniNe1T/Pv+pRSOZNAIbOMvwMKcU06elg2u/mS3DnpeZkzzwEIismKilyYYc+q/eR6dZgcyykg3
cZxc0xX9veDSC1/xsf+ODDbPfVFhf3SGFn7jkHFhGHnYr81Vnr+FdNmdVPXXsHcMYIWsEJOuXaQ0
m7Bbh1x7AYVecja+6NNaZrUn33PlLeYq36uRssLYco3UYvVCyE2Dm3nWgQXfplSUphAZtc8lhSXm
rnbsrsKvUqKtP6FIdyHgYPfh+sRlIQmYoVNanTca6WokOhGXtkZg6HFPFEIRqu5bBR3HkrZu4+De
LGLaXv01fDMAoiDk6vBsTwbG6rO5FuXewidzUqebTM+RhPEdzW5bfHyRm67hf+iF+HvyQlOJC2Jx
o5/O/Wkt493XK2JJFoqG54OWvsJVh6U5fu3gkKCqhHi4uD7Y0NjpofQsvRVmcGl+zqklNKSLodJQ
AUr/1J9PuOZP5Udd2zo/mo19X61K0XC+Vi/6/5rsMUnn69fNizUr2m1Q14G7ol2KozzLSnEoeRQ+
fU19gCWspxKnt4H9E/r3T02/7FUN0U9FGSRJ1QGDDsDXri/xkG5luVva/9AzdkH1mmfMIL5/fEpV
7jEEJKgVIYokewCCSqNLrCG0FipNmi/b/034JQgj/HWojbfwWLBZhMn11GrCGFgQCsy+70kkoOTA
8d0FZlFiD10p9OQDGB54mmE+BiuqzBqFOmKczRzuXsM5artyMkHIbWKJfDb1ixGpOwihucy+o7lA
ZuWDN2IxLQ8jLwCQeBVm+490wE/ZN1arPZlRBDkz9mk9ErX7GCFFn2hChdeqUdbr35F1uEGXUI4G
1kScYZST82WQm8VAtTRvE0xLYuRj3u868cCeIOX8+EJcmUo/tpbTFJ8SuCBqgUeBJw/6p3B67Uns
wvpJurSRp2w7fkh9DCANUVem9Vg3h0n8XaETMImtyjZwkfXuKRDsyDcTdsSBdQ9aavuNp99EqBWT
sCiZan4oqdC+BvfOZf+zGpCzb6wA3j/wMv+FTS5ah4DpHq2JH9kWHrDvlrByInii+Fuw8ti1j0v0
GqZFn2YBDTIZOYO1CKP1aYVMmPhG7yz43hIpfph5JxBQWNRsXRLMrzLhr2ddX8uQaE7Zn2LJ0Rdh
DgsjdHMLWr9CX29Zd6sWjO0kCNvQ20R+KP15QU7UiywlORbOSUAOAYeKxEpxV9FOtgjO1GZJ4Hur
BmKlkwZuAH9Tt83yHFdGRyVmFE80BZvtbwD0qEtv8PHruA+4fdoN/WXy6w01DB4ycVRear20xQHt
x361Z/k2Grvea2peqyXaQIS7cG7uyq9f8G/xy/c5VP3Lql5EY4XOcODmFjqIr+QAf9LAc2bSp1Qv
fmRm8RYfygv3bZ+BQQZloKTnylhSGA4Llyxseugr4zEttLzvIFhP1H00I/8zCXfGKXmC/lclDg9a
1LUi78Qj3tzzEieX5cx0jDjZJ9tWae5cP5noOQa6rz0jp6kK5smbsF9kL5sy4Qtl7AyJgVq+ZrYs
CKJbKoqQ62WAyNECTm60J8PHCZ6Mn2JISNU0yJMMSCpDLR8M3xHYTlu0Ia+f4H7XsqRcZmJ0v0Ff
bJJSfttcGGvUxLH/rPWn3X3XJI+59jGOYvtDs3f1CrQw+GPWSMZ0QKzBIR3NIbhQPbIjSf18GMM2
KXk4WImxd/Cqm3CjGNIj5ZoO3yj6M2dKYMg2LIahrpofmm8M/E4/GYJcp2KbYvBvNpQp/anzmuF/
4eAwvm8GHT5kJifNNd7jEo6L7QaEyU4KwtXM3INzQax32xtGyUVovLO3cztfr0WURXASpgeU5Hxv
aSE0mqZUO38UKknMAW5iyBVomtj/FkpJS8GpywHZjHmPLKjIi1qO3q8JJx0f48OFlDXsQ3aGcLsI
YXEveZMGeMMjOyteNKrtPGGGvQeNFayyutPS2rUCJ0Q/1+hic/YzDEvItMMBvhEmeCAvQEUew2cb
Jaa1QMGrmawaYoun2p9eDhRFrt5kC+vfyKsBzVHsbgQHamWc8vnWxRxZE1MeMgiVlc5MHEQnwTC/
WMp86VLIAGlEQKfbC8ZZIQtvgw/V+k8k9MTsAwA5Adx/up9aNxMajlqxF6MIvLeQmfXX6EgOE8zQ
k9To2c9QMu6aOetmud5YiSIlt6uvYdCKBny2Zq2PlgksNLhQoWoal9jYESPq6TNQMBNCcVJYJA99
zKHWb7Jv+elY1CBUZdkMoy91aW3v/9iubOG0p9Q2z/edhl6AkjnqG8qjZurJ8dJcIdO97smBEZVn
UiMfmc60jQPZQpRp8J2W/KMAUj6UePmgjG30vRHh920p7lTHHhy58sXhxmb+vH/9S7JbEOpdthun
U8AuydybkBUbqX+eX4Hv44zeEkf7S2MQO5rizi0FH3+2hGC1ML87XjPCaGFp65c6dTra19w3xEbP
wmRJZWn249V2rXjGbyNoqcrp178skO7fRJIwAmBe2CugIb1vBuB4qkolgKuGI+TaCtLXkgThhyTi
WHU2gsw5XBXLXHNTuzf6apYXKMqIMQbIqiOK+FxII06Hg0YFg6sP+OrfYaT7HX6vmfU24vccWJrS
K2U8I6Jw63r957K4V1uu/luooQfP2g0UjvrcvMGO3WX+iwaZnBSUWBlFET5I3ma7Zmn1mpJUabk4
MvAjZKPlfNm2MJfAHypmK2yKcTj3jwts8UhcZN4ylPTNOjj2+T3hfSRQbHxmpSL3DlIAKxAHnQLP
qq8a1+ZOPKW91jgRe+lC9Rc4SRsqjm5rtxEmK2Ig34GcKnb788qqBFSW5mJWnp4j3obvETchScM7
YpkyoWwjM9UcO3/HJxpBcd1yslGAx/Io6348GDnbhxXzEOpQ7gUtl3MrZ/DmnLSnhBXIZ6DSKtem
OAE2R3hLVUSTd+9+Ie1FqZXE+tLsYuNsFeZ5/Y3Pi9/h3c2w9Pts+Cu464BBPe4suYxGA/2GE138
I9ge5jDsQ6VMgpsmKZ0PkvWrSrrzl7L51J/lfEv/d9wFioqlnHlM/CMW36+w2uIepT/veIFlYBL9
jVdgjeN0ueYRduKJLOsW9rc9XlTb11P5H5EUhdhE6h8g8HaNlIo/XgfDhP70sdy4fXqSwvzUHHON
4EYua8cWunl2rWDGRmhcx8m3x8Wjz4gz+oHIMmflObhkKrD2PXNRvumazA5iNgJmlvc1N8mCq3H2
N3nn0V88R/T3D/ZgOvWupWUPQSxQIlcu+d/ctbnSFnX/0TByhvS9Mu6QS6Ger0/zMhbicC9m1GAY
8TWgwTjWV2geS+JRsbl2l0ccOuaIjD3v85jywq0Nk+5EVI2pX+fub5CFrny1UYSYAKvxnYB7rNc5
vxYNj4IKsOW7CRy7UOZK2gvY/4sS146m2nhJ5G7jI63+oN7yb7tl+gDXYHa8o1j6c7wpUlSUKb39
k3lYtGnquizsK4me52Sh/dEcJrOeGunqHuzwQE/BcCJCMoU6Xa6RKkBqqitGpAV//bH7QLK3igdp
w0gWCwQFxVtLSVBZCfa20hDDwzPJQUYKIiHJiaU7EzFXlva/WBH9kbejPGR+Tqvk/TcXBS5duJKs
zPB+P8HiG26edl04LBExzh1t9PvC6XpfeOBY0C5wUwo7n8EyJ15TtE4zYAycY/GpiX27f7qbNEcZ
ISURVIXYQQ20j3/EcDQNXKV3RQGruxQjLWuB89A3lgY2naqKO57F4LXo34KDtCwqyfIB7vpOWq9r
csAIZKcpNV/kCdSOKRN/A5VBaO8+FTbaFgfhaF+f9anLxaeF0JnAGyqlHU0rLsTDiWQ1E4ApeR4M
eHPHFIMm4hTj1nISHwFmAssQ0ULH71qndEAcMRkpOfDk3zvxAr0JFaeLNCOzwRweW5kl8NdAgaaE
6RY26mCLTTR2ddQ6Ha4Snwu40uZw7PdCo1+xxbWId4RUrQPZaAwt2+gFyJ2t2ItoEQiusqNGQ+ZA
QaGn+AomrnM0xB9Ft42hSGMZNeu9G3OBilUIeUzEnVReEde0MfC8aW8moCr9nN1fllM70LSS52Zy
/1nAh345Gqd/m/S42L+/T9aQVSXzE5vE5ykXJQ2WE/gou6BxU1VlDfT72mwhzKui01TCBY2gzSHS
k3oMyUBr6//M3M+4hgMMdMxloZF2jpXh2Fk1JxfMTR9A8GMzT/JAgQXvGUoBPMfBrKW7Myfd/mtg
RueTppBUlNPLdteSsjXN3k7TYVqprgCL4klmP2gguUhqODS4t4dQDCb0cs7n1Y6f7YR2ScjQXh/e
wtK4sifaUS7ncB6KvlKAFztmxJ3FRnlCS3o7cQ439XGlQrsjpr0diL5LcScfF8edkPTqgeh24c4M
lIsYvOO9fj/nBJvpkdShQbrNAMMZgVAsU1mAw4WD4/lI6fnFxQH3hu8ZzZiQ84JYa/QX/flkja7o
dygDITrzjHp9S1dyMITSh9WbOT6iJgZUYTFNEJ5MI0Cr/mSghKDNhqViQS+Ozn5VKBBSW+V1/rXF
bgurn75nfhe2fHlVAJ6NdT07BtD9LXP9NLZMWkz/WOPFm/CPQlKky5wmLcqnkVtSCtRO9uGPl00X
h9sKkQFLFztiuTUTm4PZyVkfK5X7jRBbDA0utUImr6Q4tlmOVPB6KKqoMg8xqxPEnFItc2ghUHY+
TsMQFTB7mNESxi9trS5zT4E2hTrtNiE5iziVlRPFB8UqKyhsLEovpSD+IWb8D817hmiJgQx+/ANl
RLeoml/BneV1wyFNrlqczryMzw/E45nddTPZQgVySrIV2vOcJmGtKNExyjI1dUKW5j0g1XhEJI0Z
UCdUsCUBlSBEFTLkJ7MTwHkt/xBf3+6aAdpDZySKlwPD6u73kv9HmP7Z8+oJ6LmbcD8VZGFNKns6
T21ty0ApCTEG6sX+AymPrQhVFG9KS7PPi8aKXaF/U5/kw6V5lJYUpSnSMZkhDI9QYtnn/s5O2cTe
O6/ZZ+jyAnl333TxhJF5qGBsC2JICYwQ21Yp1QiqAcBRuBrzBEo9zQtUR3W0JtufZs+wlgGMVMjT
aPIjsgC3xDjQfeemCPzVjZx4Lo4Xds5ym/XhAEnioCE+xQtDB3rHRAkRt4NO6gfDMJdhbF9fl1Cz
Dt5lMHK30dQdT/NIm4eJAJKOCXhMzupLMj62WEVI7rHW9LGyMcNk9hASP+JmVOELLqKiC8BlOEgA
vpigkupeCvwnRcfb+KJdwSHOmE0GN1vSjIuKqWfxSvaTmdq6ivkxuAQl5T6VR6oVeY2RXuqoW89c
BceIJbWWrd/ztYZil3P6UwmC7o9V6AnK+ub0o/AU3ZZzYLdbEAwU6BMMyNn94SJCrBaFLjBWJtNL
bI/QYT+W6LzP6OnPdDxtyXiXPZ5CbkNGQA9AM9RHxtK9Gazs8SWj2WGp7rk7xOusmwGke0xfmspx
Hhy0S3d7ZE7CfdPym1XeqToPQv3I9ssgSmyIsz3KtN79QRQM1w6P+xOOu+xcy7eSFpIQkibxLNUG
RJFGYKwDMkMxtu+ip4WUSKIZfyvKlYLwXYLrgjNt4PcYqS9rJz6ywcE1w+aBMxkytFdvg7ZMczyo
GCpgl/FWxNNahTb7LEsxmcuKnDRfT9uhatxkBarpnlNGs1OCy7r1H6OrzSHVSlHX1w71Q3meb77O
r+Zuj9XsvNhB/tVUFltuRDYVkZHBjA8LtbTMXgYKI/cw2iJyU9/Dn2ojSpoWla+5A+W6HQonfyVQ
RjEoS7wlKdmKmXYWabhKgiabTYPVEb3+okfohr8TrxWWthJu2V/s+q2a0yMxNzNCxiQCpZKf4Ev4
Hy6XD0nQbJlaWAJPrmSdtbW8ARxDe2RVEGh/BVHg5iV0qKHcLR6S560scUcrcQapP0nSOTOBa1u+
nwEXiSZgNMvHZS8/ezhMfGOmj8vz0IIiCOxOQVlGxmJQmq2ua89TRfMYOX7ja9adPyhTLZnGbgMP
vCDv3f6yY6eoZDN5On9+V4vl0ygcvkVF7fKCs3npcpbBz1zPJkyM3roADOuVHxQv6QzXwdDZYx3O
pL8gKSREKC6dxQ7OmKhNqCkp0q5Z2JLEsgEDNGK9ESUcL5P/XbrRmaerTN+YKCyXljRtNHOHwftb
QsiXdpUTb51M6sAMppzpdLcRNFtVWLim4VRR4+h7GfgLn2pepYfr9j2ftOlNtk+HeYDc42YiPe7C
fPbimaXp5KO+BPSstfSZ1/WoK7qr/I2LJqFZ3NMaopUe/CF2G2TCpVjeTV1ufd/0TcU2CzdwYv4/
nELvsUcgA/C+VoE6UjIIPcQZzl7A/PmfxpnlcIa3b8yeWWo692DJFekI2AyiCF3bY80QnTdbIO16
KyATdQ+yOsSKMOokMFi1qYVeuLcyC4FYVX64gB5DT4f9XT1CqeFx6G254XTTl6nzLms3Djqe1EXM
/ft34uIiqTx6VwQPf0MBAdnffDfyKtgev5M1YRMeYiG161xlkqgX3p6ke5KjrdZ36JInEmbOHUKd
WummqcbMoSwybaI8OfsMCeozRkQzPliNu0Q77JzwgQW+qNDK8FJvj2wqcG/9isQUA1udECqRaiZK
TkgrgHYrE8S4L/qbhLd+IwE59i+D8d6p4ZDRw8ejgseNhqMrUOep4/dMo+nm40SULoGdkOHZCVdm
xKw/yy1bkkkiEPQMRXFdq1HkuI0C7WXUJHiFCz8w+utSoJMVZQaDOWoT9rFxezi+pkHggyClyJQ0
JC/TL54pXckO7bmbBqMaOV23aaYlLCePqDVbSCb29Sygo4UHm/lbsmC7yoVHT7445MwUj98n4+ad
Ba4X0pzahgTGqc/NhSJjXisrXeBZVRCZRBfcbdC+ID47GWlPjSifFo9shKO/NX/x7PPu8ztZhAx2
uJhNBae8vxmr/rAFN2g3cAHSKSmaAQMA5v4SKdqRah9JZvWmX9pJL0zlm9bjYHSIil8CjkZYzkmz
feiEq6J87rGR7B8iAl9eFk+Nsy9sRBJn0HphyMneZj7kYwxdy+8G7XbNm+KB1UhRJKYv7iMyFOVO
f03sMY5HDvsJvMfu2OXz1smlaNdB3Y3hiP2jWjf3yVsl1x4+weByPU4X0Ix1b0zDw0Bi1xzJ/wbA
P+Ess2T3BkPZ1jGWUBmgjrHIkJfRt1QnRVUZ61GM3m5iGLqU9g5JOesrMiw/hKZcokiYu7Z0+JMy
SH9XZOlzNCIVoTshbeI9I4ksyk9XW/sKZCwbBPfOVxY5fkBj2LmPuPAy6LqKxskAwsm+17dLNu1t
ljunh2voraYGJ61YeQ6bvsVzx3Kjhm6rmiake5w/CGJQPLKJ6BR/tycZevJF17YHSslXRG11nSYQ
XN0D4emRrSpfun/bjB5P29yTLpK/zNADRECP6t5Sx6Xf8tFEXWdDk5QoaVvwXfH/LnLoqE34ikVw
14Es81CNyekXQs97dgE48pVbaAQvd0p0jHQfy7T1LitvPCbVZfhSBBS49oa0J598X2QrHpbwL++U
gUAsI5hehjx2t+0hhjU3vHxuFMpqQC5hDf9stNa96fGxWN4e7C8FstAHsecp0WngqGeJLZwhGXeQ
lPygBik3jKP4CqiVdb2hHi1wxdkAaYUUmtoE8Rp0IbXERDxvbhqPRscrgTtF3srAbUWtFm9zbfls
W91n2XE6lSzwA0HtpdPlxFS6HVaOwowsct9+weHwsaWxSKvpfMH7987OF3mra3QpcaR7NF2bz4dz
FhJzrVzMCiKYw/cGX60y9AFbTi+M3XA31hY1XmD0qpoqphBl3d+/yhxJJHYwWjSvfUYsy0b6I1RT
pz6ybCT6AKb3hEugn7au9GcdCWMyaH73OtY3Bl44iXFE5nozMhTTOuYHr+26ccSal7Cfv5QDpmbP
U5xthUG6RrLz7v7b7U7JyBoovvpCN1WN+GUoHLaoX2zHhmqX4JIj4vgf8K4tbEfcmesvIiJIyXwf
BZwQxBYSTauRJnWKwC3JM33NWSggx11XEscuZqgUQtZdeQFC6VmtOP2xSPf8EJFpOCwT25wa1nXK
Sj8gMk1tnxGzPWh5S/f4EdAcsg1iscnoEcw0m7HHoPDs2GDaAgDpTaPhUCj2txG52KGfhOg54SXv
rkUDPeYx3DJxz5GJz4/T2VzgJAWwXcsW99RLJGxjso3VFuCosB8TmYg6+5QZ0iEFIluGsic4nOpP
oR1n0lZATRcvJj0wA5BSL2zjkU/+kTb/0qmA2spO5xA/D8amMql9mmENWE7NmP+UwREmzxhAFvn3
erW+bHDZc9YXz4QbE3htMjQ4oO1Gq235UGYM4Qokz8arCms2/M1BUt741bWrUGcyPFAzIroAVJHE
2sv1QfhS3yMq7JTB+U38EEDyXPRJh+xMaxnWcwYXx2PkNNjFuHdV067P5IvL1QbFvs/HUqXmj9hO
7E4ay4sK+Y2cUaVoCVURIt4rnTrOFffuUEWOV1wgeQrpzxzaEV2AU3xaBcIOOK2sa/+D8nYOIB/M
P0zs8Pm/Qe9PeJBupnox7nBqctsOYPoxZ1GjtLeIsAIeyLxk9kiijHBlDmCtNQULHBDStxjwtcW6
SRR5bNIsvjAGiFpHGYGSvH4OcaiIBR2fqOF9crzc1V+G/UIFHnL49sAG21kdNgeqUHWIv4OBEtHR
ik2R6dtQCibbBqFfdLU4oJaSWPVwU9DD++ShZXCIEMdj83hmVK1KbljsEToAVHCnK0kCVr/X5Zex
0tpBLyoUJiegwQTZlB7wHG3NRelcPOUMVA7NJNbcrWi8MGCmsDOEpQINu5f5XndJ180pw+PXyjwm
PR8zwvd+KSoNzNiyANuPukdJ9PgNehTAtuC7pH1VGBRdYdN3DUaHCUMucGVwn+oladtudzX6HDmx
Pc7QKOJZTFXA0a/liRzhRL2O57qysrFR1bvG/7Y5koGCoDlfC2+7gdPn1SwHufKBdDpfF2KANu81
aicV4493MogOH+fvXFpd479VwPKNNCLwRcAQQcgvwWCYDzCRjXhSX8uLfcDqOVvt16ECz3tMxgIP
4Xga23puB+0qR7pHZtzL94umisXiVKCMOjB2wtXHlo00+93TrhsA7acS3dQ/Omyop/ZIBnsWEg6i
b+g5deyJeqmPHhn7rSEmZku3p40CCPDbf/V6D6hC4mLcws5lAX9EAHI3DTpWF6NVweUMVJ+D3YKd
URCn0sunU6aOjRpfV4I/K5AD1/zuxk4BoJnEWjfObDzxm7YJJIJ3spmsEdgG30biUyRYzIXJ+6ub
NntPZb8lXzOUhbQbR5bychLnswup7kNkQoOJUZcND5rP2Z6sHzr69Ght7NMy321omymTyc6/DeC0
g3VnyG89RwrmT0edcPJZInTfg0wIj5Eqw5UO/M1eiIRPv9IuiFy4KD6UHzHnebaWe1Z7Ufl+ugKD
195NwlFdAs0VxGAJG7P2zoZ17ldPjoXwqLxvBRJGDqfBVuCttW7LFUNadZpC3KCDMpMGphoc8Q0C
IpTmgLVNdNTYIcoQAY30CwpK2XPdIPpdPGw2Jbi8Pvzjx9/mUcvEMErSuqqjZThzNmSpdP0/hsA3
5PrRT5i/E4ah65gpQNav/DEJu+a2OVi/t+AUlKwD3sO9qLIAjYWFlE5GC3peemvdzwZ967p7VBw2
4NevBt2jllJk9pjywwMFEKPJ4OG1/zeDy3wvTq/J2ZWhKwXHMPnADTutBORp4WApEtW1lD145oYV
5taoKMq9h8UjWjxF1EUVxsXwRTvEb1u9ar5Bv+4pe6zSeCTrvcJ1e1BHWj9VBjca4s1C7fYZvt9i
K2nJ5cuHge6rR8fu0DZKGX0tnvDD9Fm6ynpX4sPjsvpK6BmmUnJz12uuvyZwUglckS/Lu4j+DPE0
Pz7hwU8usy1+6BYr96BgX8A80Z+/HCqAGIMI5kIsMJDDhNK/96fJmxTXYWSIqTZQITOBglY3WSKB
K7XDYS/Zrcnq9wEpn1Km4wzXtJILbulgeEuuXosdUWKz+7+VDtQG1bnoWpOuW2W+TccNaeJLSbcJ
e1CWhG4fjgSdHmHzyA9cQ55OVldG7a60iRbAtRk3W66ljsYsjVWARORknBYpYOKR2DUnYfGOeb/Q
iLt4yMoKnUWZCmhoknmjwehGxEOcvoDF+yMyHOmVzJF1WCA2GnuSCxjyoFKBq6ecBRWVCRLE8bmo
o/vtU/wATL5QqKrLG+RTfOYEY1XOOlpb6uAuXhlYi7ES+0Ulyv3A/k5tyAP6hT8cwTBUTzPK5LjM
xMP/RIG4pwj1mdifgLVq3xfjXxQ0x+5zeOJ7nVhPiTG8UcGoiQ8ky+A6XsUyhRAMqawR863URWSk
o3lLv/4IMzSjEo2Y/Tw7XvJvqs9c5Ccm3DZ6KIick0N+CUbuYXpcmhxFTya9G33CElXS8PLQBBZj
eEUgFvTUDpPEAZwLJ6wadRJh4c7BDCsxIBOnpDzuCtSofnfaLqf9ZE2UPpuKCtXj1VEwZVfdrvIb
GA+Qwx1KoOBSMz2J29g1xBIEUxTZMIEzaW/Vd3iFFLExvTodBWxlLfdXIm4B19IJZyBdctdX+XTq
9gtk2Gfae1MkRJ0hgjyhDF6/Odu7encSnPiZpove0xf6rdSU2SU4JfIg1ZwnkG+KkaXbh/81JN0/
/hpaCBq1+8qtiGHswTB8Cm6hKip3jfMkZSzCZg8atNt5PbluGzedjVJlVghYfdiNkXLdnLOATNqU
pQwXMROIKBE17vrfQ1mvjrSUj8c2bKgprxyxL4FNm1IBR27Ead8e/9wZ0UccyxYx+XvxR/bI7NRm
52LvhyghVvJHyDGfvtNz5rk6PSHnE8fZL87ChDXtdcVdPl5FyEQ1yNdBuK55sdEL4xP+Ytr2TM41
k3jgqXcBS15EdY9cLIkOo1zDKJrX5TXDZJeqXIOceKPOx4u1pdafvVcHp3mbyBVWxAc8b8SHo3bc
4Ct/GWXdbkfeFQOe39R0IbKmogjN4QJEK1pwjzLQ68FGlrgGjxfsKXaQKkr7wLaKwN2+VtEkF8q8
tydLqrsLWHWBsTuxhiU95Mw5pYd0FbQ5pbcZRURvJXqQkKTXXjkPsYRyAdsrWFuTkP6V7wHh2DDM
58mJY8g+us6G4cOWi7hBxKPXRnDIULwe6Yf4LvVDXUUda93IWZ3VW6tqq2Bv1WBAmXMVuR3osNKv
lSXGqkWBx3yvuFV535kai7LvbD6yAHD2jwtxsXQRv4qAdwBEffQ/gOWJtx1X3ArzddRZ9O2sk+XK
s4H7EV8VajgvsaA3XUWH8yJZ2oaX0i6thRmeF+9lbTbsAV70s8AF3orNSrUcMMiOyz/IHYH7Gp0X
ld8yf4h+kEV2Ko2teQPZE/u2JTgu96Wxk9c2DP73LCq74Uql1m5DUQ78XGaYCA3ujN8x5qyiTtK0
WYZD1fli3wXAkgbzp5th6ISHdxBNqvJyQZNi18pV7dLq++5f1z+64lMNKBYtFLYVJc898Aus/2lW
gr3viCaishhJdEWcFpf86vVbn3JigFOiZC7mnAIZwj092mRTbVOkVOoVY/lv9wWKNtWAijzjaZSZ
XZriJiPnyypwXbQW8hIZ5HGtlRnF4sJn12x/WbPKX2DFGjKb2Rkb0qdJsq8fYJJD22N3P+sI0j8L
oLeUeJfCA1Q7+Dknq/ZPs+xVSlIsfA+sCaSug17Vov0tAv328wSQtgrZ6IIrPGU3QR8D5pvv2Knp
R1G1kPknGaOTnCmJOrbTcWCM5Ox4sRsImnWX/yC6OKfyoQ3m82pUSSJElmXOKSw3ye/Yi0qCduV0
b2xGzmMXQ2cj6QO/PyiR/2TlbeJ6g0AKfvhElQKJ4kPF9hncvxdQTksS7hl0lBiRalsvVVeirvy0
eFZiFMwiUH4Fcasw++N56I7StskrGIp40SmhzQKyp+cHOgGweOW5AunsGhQG++pTcuHPfIIUhZMM
O7QkuYXorCVTuZQgnmhd/WL2G6FhuE+GQwSgeFBNPm+kQFxGQV0Xuhlj8F5Iy7+j5B90yHTQXRIM
9EbjH7IfKQz+lg4JeuDBIexpbW6ET9izF9TOdEbbRvw4tgWzzEKG24E6mYgTm5flFntWm7rxtQF/
5zFNd+s8pGhhDlH99iIX55Vro6rZshUkO7WTL7CQre5v/QZismaX8hGE/ai3dUcR/SD1hu5gEquj
MmdBPBX/Wd+OIt9mF0PQN4d6P4C5TkZuqMo2TXVLe1wTGHX+jBaZChtEb4iuEgiCEVhd941MEFdv
BCZU2G7FmM1Xa+UI2377+N+k0HAhGnGypwZDN234DjQ5tYSE6MV0hdIHL8C3xjjLkOwAZ+TaNsxR
Hr03v8JfqyAmUeiooAKk5Pdx49bxMV0htfIMoFZi9DqieSriXQQt3AcLu0TqS/SYN6E4MTqOI43b
10y2ipSmIYmeZdzvXw40cHGUujjKKcNRyNmFcucEwoeXvbpaYyDvU4T2/DFpRyUvnSxjX7gUpImO
FCuOZd9YBxKCWUtzRJbgxL/9OpY3s0l3HTLhSF2XTxZlnWbXZCMBlaFIfpgG9OXHQiCyjpya15oi
44Ly7VR4FsBZkEytO7ebMKH//qw9u5/YOscHiArWw9u+7DB4CnJJl0WhBiGkUNeE21lBE1IJAlZW
5g3dtFqpZ6WIDHmhukmphpYWKLeiPTNVOeMBqOYQOh+E7sZ12mR2p14xKeWKfoRUSbg840eB7In7
8Dh+lktjbJLJjBiXxlY9zTMAqRV0RJndOkYiZU194eoaIDrGSV0juynfVWJFaeKQX9GvQG0UQak1
2+O+qRKoKITroQZLErJZ5skzxOfxBzUzNwtG8ZU8nA3NyvtxNLp35PLJ1dRhjBRG5zM2DY8ZpDA6
VYULibufn0MsvqfoP/YjMEbE1DiMwZG76kkE4ZaKI3gkLlUHkQuNiXN+6r00LsuEhb4e+VGeeRX/
9qVOQDn3mxuh7dCpFbij3Nn0HFDblIU/0EZgXYt2M6WBdt7JQNBEbz2RyQn9svwhgm9he7PlhZwV
lS0j7KRYDEnKU+kk4qtE2pzw9UUj7p3T9siYttqnDVjA/KGPQ0R2rccgccuUwndgE5ag0MdoYrTW
oiM6lyn1UcTdVfh2SBTHY/eGWHr+CDa6Fp40fZhIpmCJfrJNJT/YwKmuwcgO+NU2Mj/ds5AT/biS
HBbcdUgc2mjtVgs0OuXMASunZT87kMSDM99O1OOyyeBotxq22LusFwQ4NF/BHsMMDjlZ+Vj4hrLr
5v/wA+mByjWuGcPuRhHbuM1xirxo7ty5daVAH5T/aaOs9GfwTpratb3JldO+zejd417lwlMf11JF
oBQUmfelR1Vs/YLSaaI0QS5oMvlH3mNvWG68RjZdGreGeWVzgVwau2IPoO3HjNyqKs9Ve63rmnk3
i2vboEDKSyBCduPZkPY0pqywFIyfElH8TZZPEJb0HFvqEH3caAvVIhC/aqmlHKDrEzu27SHBsjIX
M9zO3mtPU8czNzd/9syKh5LeZxeOe5cDPZY4PpuqcDk47BuRoDRlRWVcehXhgOVAqmLnvOxl+SNd
jWKmyI5c2cHY1N4GrGgFe6iwRJpgy6qe8qPPAJSlDzq/YRYbIlz9IRQlOmizZpLrCcjKUlWHKZyT
GsFUfWcYagB4qXes/N5uuQXOKtjHyAYKrJ1TndFhykUgaZw4wBWDZG4ZoFEscrQ4Gejk9tX0Qmi7
uwTnj4+X7wPwztzRpTQ2YbqRuM93ilsMtDRyxyOKjs8gBJGYs+b/que6mYS8Kr3uQINOMVI0dPtS
fJySn6wmYm0Aan9vNFNBwoJm0GXPjtalus7lCEiwTf0ziNTlqFHivYzJKodk94zlF9JNoq6A/+vx
bSJreQI9oQLFHNHsrygU9T1uZOmeCoxrcmIeXeY0HC/0Xpxn6RefoCbXLfGqwTwAPzpX0diiRsPS
hTuOMMj7C5GaZiy03qL0iRUf1sPFAp6XEb8oB7i7MOCtQoHECcvAgM/BKnDwdYF/Ul01Srt2Ki1k
7mMeZyMuY0hsajigAvFh8n22Z6VQxHlhZeasCzn701BqR+cInMBRaubzNX4BcNf5i4+lroyXarpx
gGS6IVhdTQIbzAn9WXrEXqjop9pWNsHQiY6OaHbTBHm+rXxV7ru1PemdA185NIEx4oe1/MInoKAg
UKrqtX4MsLL/Yk+RV4xDFiKPkdagvpkRv5vggKdTJ3v+faOFcKneBOCn2CxutO4BWLLmt70jwDFc
ONqdHp/2wsZq4Ghwn41+414Ci1srSkHzSMpPh0IgxwlvFA+0zuGsZkUxXrD36U5OJT9Oo2BaXKeE
cxc2AeliFWf3FGDaf7U+Tvyf04aC++/hTixVGjPXKXar8EnxJ6ZEZKywwUkxK6OoW1GlImB0eE0n
jitHdcHt4opFnn2Oo6yeNQQP75q/Ha3jHfUooIEJLnNjjeqc/WKpIK+ID1s5LNvq5vqr/Wl81Soh
3q7elRwiWcpRf1Cyx/gDPRkmubjhH/oYIY8s0ywGoM9S9pchpe1na3rX1B8+C62Po9vHVBcz0c6S
toM4S5L5EovSFWO79ULfqFH1fRUUCIY3qo5kWQj5BYsczaiJTBFcPc3CW+u4jiwcTdmL0/XlV7Jm
sbei8ArUwJnA0SMXGc8naRcep1d6pz69Q6xvyrnONFi1qN/8nM7hKRRUmeF+veliOKkCwa2Bjwzu
Kv7l2kSW4sSISS0fGV2P64YCiPhsKWlqPDP+b0e393UUygsnKtGtVBJVaK1UAbNjqr+MNkgSuWhj
0J7gwV0dusdN9pEMygMH6fd3ffwSwMrwucQ0HKghhn72fzhUEdPCTmU6yTE/EtIGnZ7DshzupftH
/tepijVwCzoWR84srEUJVvVqKwqmxsp/+/iBcEF1WY9Ijt+XFQwpEEiOydf5OCDCr4xfeJG/q4nO
s2eTIc0mkU392Mv55WHdJA8+x+ArUdhTaSTznWwZ6dvPkmGKhH4ktU254d0fRTBj0zeYNNWfef6q
A64ExOym18OoNTnbD2mRGMLeGq35m5pqK+ii2pT09zoFWjs67gyQC0DBsPAHagbY23zjhjBlHMA4
WpFwJNAWL9uTSo6UIw9CyAZ6XqMhXKZOE1Qa0xiBmnSacYsQH3yvxfh7Qb84MIklz4495rFpC9+P
qei2+es7F7O5qMIIClEn1vTwexNs8W8BBmge92fDADeMwkRWoCvxWTKNJcdlcHux0HjFhfupy2zB
4Waxcn28f9b2zbJaGYzXzS0ZWvYruxXpKVoD4LXjoEeXdQ2W1fTf4HitAc5asMp2OlxG/gXZtO/3
Eh3Z9TSoLpiuPgYa5hwULi55n+1+0y7MNwxWN4fc0bW9RTGTIGKr0u7uu78JkYsGqWG6sZ4HUijP
u5pmhtJNDHU33BqnFEj6GBHajiIbMiBQGWrMISxp8mlBCS2hfI4TRwEAcVaRqSM9hOtRmxcYCLKb
PLsHYVo1Pc11zeMhtf0fpgPg/bLxcnTNuolNlxpPH71k0vMElx30GMymWzQfdszFYbK1Su/qUG1Y
5NLAPE9d/sG2IIhiySRcZ8Qmh5Y+JMU9X3bvTZ5ToQZgq0lo3XTeHKzKbNtDt97n+oQtw+F0mc1l
LPqod4TFbhlti1LiKKRw6SdDEEfb72EMQTaLeoMLedP1xEvM381/mmI1HBNUFTRTxuBDWAnVJc6P
wtzazAzSRn37FztcQfTR1iqHWeI+o4CXPtGpminsMGd791+ZYKLVdttN1ruXZOjgrWJyE4vcg8H7
3ayFFF755Kz4XO0uq+oj4Ge1VZgrrEtnzTN/iauhDcGqPYUW/zmADdIC9pkBDGiUlAvw9efNNsU1
GaM6eo/jLeGC1kiTS6dN7BnrwVp2yd06dg3rkCaBLuutCKRbgFp3gP4jATlwWdnic4MO2qHcgj+h
10ENdeio+0KrOZyITM8izJLC4S89wkbZ80mVQouHoGtB0wqKbQMVsJXxtjGD/QOXXaM1eoG0gWpM
KUIe3zIBQpqB1S5rjuT6Y9McJxugcK5Hxyox/pHUpXehsdPKucuuZmsB+YYx2c/Z8S69s7d9LuSq
KbpCNo70/8U870Ac/fuvRS3uKGUsXOT4tWnFZlmFfxEGrZPWoDhSkjM56iseRX+QAMeqJ6sOUeGD
Zw0V3U/LUxjSP4Cs46TRl2YBeNggF4XTtDc8amtpBb8VQXelm5F4U0RDVq/mP0LzGLgtPJtMbGpA
giq4J9knKoz21R1cxww0eJJefpQQKe3zfWra/MUiFkn3ZuyPcHoli6bU7Y0FhXM4xhlZMSCXYCEa
QooKGTOsDt2ca6Bxgbx9FAvS8QtxTLGU6PNfaOxVWMjIQNVdR0fgavgOhvY7xiDp0Na8Pfqs7j3n
IQ3raqRm3KPmJnLc/bPR/9jDmdPbGarWBSiwkqqajL5IyUYc5HnXw1YDit0KbtPbWhxdSFKUOtgT
KRwx1j9H5m/92jbKFBUy/jjrIw+3EmSwMSf/b0j5LDwlFh/nIstJqpIGNhlIBv2VgRQXoCJsbGRY
o3uQ5I+ZMD0Qj4RLMfqKnTZ8lKSwPArEHqs7zSikS2cqNLJIeCC2ODtTKDBBUHS2ie0Ay/3CicJS
PtKIwFl4+nvDFUOWd3uHY+TbjXSKOEBxG0iwNoNqs0MEafuIAF4iAiaV5Cn0KzbfC0s8d5ys+rLF
mgYumzTy1uOjo0n+OFYhYkEe21SLB+vLKVTZwdou+3gPgXDSv85h1lEW/JU4KPhCfmaMba+Oxosl
E2dLJ1/vArJ5Pmc/8cnPFwnggJvXTS3zJ1yllgi5fBpl6iBXP2pOQai/Ox9pXYYfSnRpgXDXlL0j
hAC445v4SElHGcfBfDQ+MhS5bznlgwY9gVajbEH5hFXEeo33EphDe/KcNMUcTblnveFh4Vs8llez
ICHK9Ayuhve/loT4PeQmxU54QdEHaaDy3FLoUnOivReNbPFK+26F/oBuL20idRgiXHIL1gcQ9GCV
UI2mKyUzQCeBa5wScbY3ukps2VtgachFUYHA/TI9MlgEdGNsDghfhuT9tfklWJBlwPiatC3UXsix
mqSj7SxBintMOeaCihRX3v46qARBDURkF4IRtGMuRgfn6e7FCgUL0DgovJX/CtA455vEheK0pG2T
eMarVgBxz5NZ33w7cI9EdDkkmn+7KYkrD1f/A/pS5q9ZdqyRarNc05BfAf2Mjn3xGO4yu8+f7ALJ
AfKrvUh6OFckYrQhSPXHbHfWBA3n+9Rjnw571yzT4dkejtGnSTaBr+02UgiK1EIKcr9i0sG6ha6M
fI6x9fdz65sfmjKQ4xHd6S2iZ2AmKqoAif5nvv+9lg8tg5M+7j411AgW6s6W4+p/zSV6PH4Y60O+
X81Q52cajpSkU3Knr3+kBK9jfIrlS69zEfoXiPrPUb0CFvfo/IhKJIKNJSYJgFq8CX8S7f+/dxE6
LIKQQaDLOqU49sjeD+TqHJsYqFi5dz5+XDXzpOktPjyYxlfDxFmnCwEQftXT8Hv72dQZOCqneUXL
hut5hDtxLv3tSPe13TqbQxv1jeZRSUzbVmRXxofcQMg6EFBMDQaBnlbM+DOkP5yAUCVz8wo8bRWB
W+WZyAOn692P8NShWjB4lCqafZzaRqSWmNg3Rqzze19GzQXIj98OUSwxb305v22SLVtc5Gbm7FyE
auGYYy3l6u3WK2pndCG/tM4UR1Z6T9yGGEOErBGlpzwRKW5PpWnEsksX3fI2aIZCPTlbN5I6rRLk
9TAoEw/f9niU12qir61kPq5tDJ5Zq7aErIo+We09dARWdm3WrSdS0d65n3OVWyxTcCe1cwBlvoc2
mIKw8Naq5bY/8wHjt7fMJXZpibwKy9j48QVxrXM3NaX4ZVj5dTnRLo68XgWqXKKAQ+tiyL/uLR2k
LOy6yphi97NVgHbfcXxRkPY+yy6CuQdSHfQ9XwBjssLDqQvXu3370wWr/JbUtIFJcqmT29nQf7aK
as8gbMY0sA+YT4uqneduRTCe8yL8eHEy6kE4zGgNkf7NqC8wmnXR9f/q5f2vwdBjFCLZzfd0IOEW
7iLt0QKDjL4WPIFN0nkPGpbK+ZR2hqPPqR2aGM8wsr5aKDxawD91JQrhPmZVCuL6l/BY0ZYeAlnW
Wbdx3HxessMDITVVTZPlak5L9ZSBfAYIa9ZDV2xgCo3N8sNu6Efj7auwkEEQVI4IKJHMvlbyYyWU
LuWZSV4kanbAhvKsCD2DS0H7dZS7/1x28x9keN9mDO54i0PL+F2oG+SVoSmcVYECMocwbZC68NL2
KefAUNC/sAAaNB0rLAzcLlpD+72i8W3SuPrLqCTt2wErOLUVrHNbhj0JbD3LVaH+yH7Mo3sKJmxj
AnUQFdrs9RppNnv4g5bYEeUqREijyiumte5dyWxnsLjSasUi6gOyJntuHGRQ9k3IRTpasHjrPbh/
sj5zYSFoB0OoJSdl0UXGJBzym1yxRxnC1SKawoB2oaYauuNJQY64alBlSZujDkrd0NBj4JBAPtmJ
oJHY9RmTdbyzaXyM2fbb+6rnq4+831FrCBisH3wLN+Y95akYuQoVhll2R2tXoS9uPOmfQQUEP0A0
Carz9GwGvGg+7LwJtod+hy4V3Ugh4+VelwMzvF+zNADSfs74dM1ljbuz4KCKAEJ9RkDs1JmxiU7K
fVUvHElwXxf4JXp2X/sx3yBgkZtiBc30gy28SoTAQjJR8Yzpey+90bHnQ6QrlHxLyye2UcQFfs2h
Bvvc2mfEjDyL2k6CRnpWfT9mOn9+FdLYjeWlzmVlLjoGOxQSBNGLwJvw6GH5MqswsjKvQTCextJ2
bYFhM89RV8DgvIKP4ZSEdadBmRGIDRKjYxVMbw7p4/013TGYMC/V/rRvT+ysDZjpXpAob1fgadlH
ej5x7x8TTjNP/o7VJmFrrNcWRYrRy8W9LH7R2riZfbToWghLXX10oYh30e2ZgWuUDSDFgenoa7CV
HZBOksab2HxlWUkgn5bzS/yZ+M80Nx8In/xEP88s7skTLY/NdDjk9z50Ilxg6RB5T2YMirfL+Mle
yuyRTp/qgFANEaQc94dl9mJ0Qnx04GYDZuqr64fuqKRGTF7G9p5pNlCyT3ImfFiQudb0o8p8JOv+
qn9ngXqWsljpLZ6zDRIzElc92xC7kHd5WScJBVyy+PYehuCpj1Ft8Tw2Ra6wJ5NiYltPV1Mib2HP
lSYee35F36xHkor8Onyzozr2QetD0hkyrbAYd82Ygn3kbHZtixTvlnudcUaHYM0XyLPFc3BxPVV4
bnbiZ7EdgwBqmM+cFNpBFPaf/Uldy4lDUFe1TvC+GRCRahgQDJSP5z+8zc9BNyzLbDz237VytrGR
r6IsqNt3JsFpkaTKyhmkGqKjlESSaJee8wkOZJKfBoB/YNXCUqC82kP6owha7NtM5t8gg/nr116E
J8g0NKfMazX1qowYN33EWf854uku+TyoalD3azw/EUzj7mbQVP+hT+lhemqbEj52uRfWsfO51jT9
/T3Dp/FxQwX5Z+x+0x1/JCzA9PO6Z07mWNPPGGIJt5b/dkTnsPFSxF707lEUNI9b46hlW9PKDqSU
r4BbZwKIdVQAILs90NDLd1JCDW4gFQM+FC5SBFyYsXPF6kpx18fJDQieEU7u0+HQARa6BNeOxBFN
VN0IVi3CXZeImvGjUB8B5Gxhvihv6YyJWU6S/QNjWT1TtIxSJu010eRmLa5e1H0oGtewVvx5cDou
G/EekNy7dAiGojQHWUzpX376cG1LPxMu/6B2hnriwYIEVNNtmw1ZsB+jOWPo1KbhKRoqX8aaRzGn
pLzIWhBwx5PLjsZ5pDuem6Mn4eH6rifKYlJqNma84Shi2IxXMvV++F3CKYFnylGIC0HF7uCzOUXi
nHd53SwJU+MaqPubNN84QIVAKbEE3dljQ6hwDFsyox/U8kjGn/pc691KNOnezmJ/HWI/3e/IIHv5
jiiNhvfDYAm7j1r5Y9mc23IhYKHL2EDpiYrqAJUjlgFwcIX+F5sOzYBsTeyZKwzaYisj+l1HBF57
LDQxy/LgWxHTz1EF+MzFvZNJxel68PC7hew+oqRPSNuTPc31+iCjzeOfCDj+c1AtN/k7qpEeAxVL
hcPwFWzw/fZMU+vwYFQlECjl3AQahkd51aheTdnkIqXI256r1sGWy41ufkIwS9Rtilc9V+8LTM+P
vhxfiZQaG6mv4pleDxV6ra63GWEN5vhKlKKiV9NvmPDkU4geYG3u3uzo7wBWcl5bhaKlqTOqhVHR
K5bU6ijI9EAeXx0vx/0b3jJPRA/qx7VKb8T0BxghCBqV3VBDzi+3/NK+e8+Rscr+ALeB/hmQh40w
1qA3mAnqNPTCnJn9Ekm5tDu1IdpYjpOfIjQH2azNG8tlNkb5jCN8y94T+3+pUxNk4Tg2zsJZWSv3
vfXXAPLnvqAeEXLH7KHtTdjJwTOPqk4RYriG+dMkN1jwOOCAi1BQXXRe7BonDpIDRX23/BTYRDRg
fVtkg0ADtw1NMDJAcnbognR/Jd7/tDcxV8P5EuK/2ICo4PVyB5P9ZC0nORvymlbWONvgW+Fq9VJB
TbesONXv/lYhAdyZ7Ys74+HQZaljEhpTDBNUCCrYGpyKVWczSvVbrgvPVWZBckDypIRasbCADNn2
j4cpnk6tR6B/tpPHgeySz9ftkWTjMYlYoWsG04eijcq0dAIcHRsfZ38+vEntoorx6rPKNN+xDVrM
WQ2Pih5xXfooMDgcvAq7ynHewPjLh5anQ9VicYCFXOXnBswjPEWfGvwKCe2WJz/Nm+JCZZD4fsWz
lRLdcpcQoJtbBB074sMBjbu0ADLRMnHZD8hiaEqo7G8i2OV8OQfjecyliV7uh/7yBPzcJjdwF7vQ
ahNll4QET/jl5hAL61yymZyYdjl9BUr0nvfvQIBBeE03aZPYF5/h2kH0WtK3e4GQhUBZeuUqAMD5
LspSH95ZAPqsqHFqkQyW10STetFtZfnzZXL4lOrNp/HjTSy/tLWMQtUcJKz6QY0m+aV7OtGobkN5
4XraSjNQ8JqspbuGZsX9JH7akNZ1dxM+4u6AlEr3HfguX5Bl9OiGY35T2kKt6dSBxu++GVKriP26
Pob/2S/0JvUzBGbCrx6D+dAQG5EkymDVQjLnfpv9t8Lht8oX7ZSZDojKzV4pfb0wCjTZgO/qqZT3
wFAC+C8gczt6mSXQgLIFgHVwK/Npe1+qJHdlrT0eKDzTekaExE7Ngz3uTZ8fswxSPKzWJwH/YC4W
EyGxstpoIpy6TW++Iv7p0GHXfjuK0ivMs9vuf23xgPDKwhdEzWBO56kheGV0jNlowkHq3apFuR5/
y9kAyPvSTb2t5S/RQin7MGXP8zIWQKKGNs7howT4fCTaDxcBIaMCTJQ49c6L7Rhe9ettitPy8Kav
9gHgnHBAM2U9EaWRU4pBkxTXR7ADlZybuhBSPRx6K8ZqoLicfoiuPQC93xsDqv3fWv8N7qc9DY5N
ZPp/nRPjEiKV8afIQkjLnvQEl5Iewt7NAa6KEisyBreKYs083IRqVNK1hBPsHeD6WaitEZQmfXID
LveK46YN0rS1ebAyirCkI8BA0h0FACJ1gTca8WQy3HGmoertMbaiPvgNlaEw8HI92v08dnqx3Xdf
AONOzwTYem54MbvsZl5ufjXFVZ93VO/2EOqPkfYbdcLGRQCPVG05L1jJDJP6ZrJuJOR1/zEk7tGR
c/fpwWrwmuir46jDyb36gN6YaKRHPW5PN9BkDobFfiT0TqBF166AL/WMi5JKV1w1egkRURDaYIrz
KxePfga2+f1Dy73tm0dS7EwYb2CVFZGofGOUbZu2fYBjcCr3sQDF4VNMPKkv7m8Q3BT9ibmawZtW
UCsA3apyMpTYhjEbWKb6LUVdVYc+BshNRJaZURbRvo6OCPbHnSgFbLUvHnYKqGRII1rIoahCc3AI
VnVX7OgfAClth1NaQkSdtTJ1x2NIt5rEIJv5k2VKpZ7HpWV1RMS/YWBBBsCB0AT7gaCjPXkqJv9y
I08CbwysVSR9YWdWSx/j7O0P0mBjgGWrP9vgDINY0WepyCGtkjHqzJAOqMa7xe/f+zqJmF4Lu+NO
AA8/CU5UirYZEpOBwjuVglmXV/9RVOV+nz4c2lkkO3r0fun2dgH2izzt7H6NnHTT4aS6L0iWe23Q
AIZ5/5NVt1g7Js8fpCyV6t8fKM5AM2Qgj+olViioJoUrhzyK7EGsDKaVQWq7Ts5z4IGQzwsBrdIp
xqUSeY9Bzx12S1EPbDp31ftvqlLgpx0mJaaxFrkUkX7Rwyl5ZXCIjRv6MNGK2NsvZoI7DivwZgD/
kWjrJ2gbKbKCiARfEWxBZL7kzjC4r9WKaRkJFRoo88SZTVAINATtz3xMYRVLmss96IM8GjDG8IZg
2q1ovtyy77tFWGXH9GFGcyPsSgCjtt+tsRMZRKJD0LWo1zAVMZAzf62fHMYx1ZOdMXd1tbZOgIdB
0LrURbnbzcTctw8P+8/+YNXRyQIxOwYKl+CKDGPnBZSWw6D+L2Zv9Hr0RFlsjb6SFNot7SIpfL0L
OjrK1oINRwEfqpKi2fHNJvIcf6hdHWUEB+H8x/2mz72WbaKyXGafJ64Ng0bQdgPLZlBDP9TVCvv5
LLzmkJA+AHAqoKkeqBMByycO5hBUY9w7bU4+9Jvz14YCBS3NugVc81y4bqj9p8MBOWajSvEVuRjY
+qiLNEQB/DfPQB+81hnIjOsele9qh9VdjLuJWlMc+RNL763R2V6nKPcMLIIpBd9hYXWxw19Zqz+0
MVBHjcc8z8BRVAEdZESglAziNEct7EsUvy/PBk5yLelFHBwl4tkFTUFGZ3qzPUPbDtZY/LCdrGHi
iqajjXX8K2Xh1/mubh1EZpEe1hunPBCs8zwRHU6s2dPBXX6O8XQBKvMvY/NSjp7ubFa/Eby2/Etr
F6DmWeXQjVBXtnHS/wJIBUfkbWMDQFwIcj4EC07OzMpPPALyIKJC9diR9PGhfGdIwdaJUTSQonbl
+uSHq6FJSJmIi1VspDPHn1PFRN0lnMqvj9ba/4LwPUpjcyhkvxZ/34a6vqClBdQP4Amvwo5ySupV
xf0icjGCJvrbv0XMkFIHX81oYbe8sYtXevVFI8M3+WdXPPw1tIQ4qxUonJpB6lpy2+EK/7shvoK7
sddIJiyZJdoQYdMRHHZHYQHhXfFlKxEsR1s5v3W9q95U1vwGLM68K5yHLGPwL6N3fTdicMUnV3fm
QFzzOeLc60aLiI0Dkbjc9z4geTsYIzgaNWNC5AOvtZzJppnbjvjTE/z7IN6bVxgBHeJCMiCAZ4TO
b4AXoo4Wk0ZB9Ie1mieobWUvZUOXkSBPaFEmfYBhiKxbPQBOiWlL0WzBECF78LeJl6QLcZ2TcJcs
NEhRQ88+stpXPki66PtB/zmh+MwhpQMbCAEi5FhU0TM4+eITdzeUUkRBsIgz/NhpYS7DgHgIW6Pe
pDIMJhMpBJlbHuklmspaR8vjhS+f0BiWaM7cEiiFyXxD41gKOYsgQX53b3mu9ZE9kJQtoKHoScam
aeRlsL/NOjfdqIhjNERw1PtysUeWoaE//ddSGyMxsBb/MHRibHgioNXjkaqoT2M8puL+T5T1FwA1
MMxYBgjuQbDn8M76w8SQGSwfWRKnEtFlwTWxo37QC9hauvak2bHXNaMR0gT3SVFWuCJGZdJe8uAb
K2LO8/r4fSLYvdWES0B0tKt2TfnebBuROIPGoxq8Xvt28KyqMtLIxFQScdMQHb3oRWemuZr8Ynmb
WGgEdCiPT5Al2QRWuYlHq2A/I3sq+i/j7Bkno/HWfBwhigFLDOf2X5bISjUXiarU99wsEXhU8wo5
h3oV/P4zzW3b2AZPOp8BWCHLG5LLc/dPd7/1Mw3FEC4+RPCuQgJ9aS5gSF4gz3ahbJ9josULjO2k
4UzVHM2QBNot2lh9Od1Hj4gIEn+WddhoXuF6DeEKEyFj1C2jBgHT/yz4yG/BJGFF6+TKUTVPRkD+
hRak4CyVzN1CqKsKLlp5742gxIWqOuqwQknbrNl75G3K2LaGshnmjc2MpV8MRwrplmvOuYH8R6gY
1RULYLbzU9cEGoNsE6PrCKTLfkUk1BgSh+NvxbFzN3WFUNttUZxf5DzJUs49zHAZPIHJDIsj0cG7
0HynLy5pybtTB4yLQSk77gw6BXAO4rWznUlI0DAh+cf5/bbUxZftcViC8X9q3yGIWH7OGb6NEIBA
nbXAiDn19HN+HlN4Okbc90cQ0bA/40XCbU+ecr5YVUSisW/rlMZKkRXUfN2zA0HpqlViFR6pq40z
ZGNa+qBe8oX04oRMUxxSXLyeqOhDDrYaiAHPxi8FIx7OIBpcUcNGsHastw/mhHb1zbKa/00SfUnz
RoBzYsCsW/xStxuxsWIEegSTQibgY8rV1/J6JDDG8+fljIXeT0OLHTM0iLUNyMwK3VtiHSibVpMo
mii09zAeHwuDaUG6tEBxU43YSkJ7O0qPfatj6WVXOQPmKuIO6RvR44kzJX1Qth3hq1CW1R+IXt1d
a641gZcNuLQmqHbyBTqcf/Rr88gQmy1QaK8/4P0XdmyrepcOfq7ZrAqA8ETgEe/fd4CZACSJqkTh
IdfvSLX+b7jZZBmdGxn8/P0Ug9Wr8IfrIX2cToCwCGxbfDKcFnqbFdpxfqbRB7geJ8V6IyvCLkUY
OUmscP34aAY/k2hrgvZs72DImioe/NpKi8ZmVfT9gcdvE+HT/pDFfZ9Y4m2N3Z8pJok+JvT2fMAS
NNbSIwBL6A+BAU3KLU4O1DjF1gZ2q+lnBOpWEKLx1s0wmDyrWYbaKNQ2w7trq3Ya/sSfOg3IeMHa
Sna9tNsx9DhT12p9RgUnUD5+HglLax70trDMWNKYSXecbR8bNH15nESBIDup4VwUghunlOXOJii0
yqF6kjUedYFrI6+Y2cBG0RfoDk28U2MBJyV1OmLMJFJaaPuy5//0T9kKBEEog6d/JMiZMuGfTS7I
uTQF+O5oC2kKT4tCr3LI4UoYdXt2kcI/Hb5zEcD6UDQfSveTGvfjDwA1VmpDGoZru+4FhFQZ6Is6
NnT0mtvPjGxhGrVhxoHF5G9kd1fBoZEEnRBOWd3YhMT3qhRGvmuduGJCf97VxogVapEPzUepABhI
UiN1mDBNM9UqtGznpNBZoLKXWKUH5SDD0AN3onXzxK+4pM59WmT5XpePrtapG9EgRZR+Rsm+4fOH
f1LtJzBVy1g5xpbGdEif4F2jBzaLD5W+gTfMa335zeBnJYJA3keEzR5weEoK+iar33Qxn7vKLp1U
Y9QdqfLPtAbPhW+uvSQyK5OAlWalmVNI0x3K82SRulE6L0ssM1Kt2pNt7lV48nqQrfcbKACPEzqP
LbNeVCCsc4F6zX+3y6JNxztL9Bk/rjl3com1wnRavtp39GdqkMs5v7ICz/Gkj57Odo6CO2aYD5pv
hIbxLt1PY/qqHesPVpq0ND3ukgWgKNVhtmggvXRjo9DicYW5JboKxlXjBfGi+ZwiIN1dK228S8Lv
/bZ4JTpTlDG5PEnDgRXxHZ1SExWwIKv11V5AzMFAg50YKtVs+kFBrJ3s3D0NHKAtuaWA50Ag7Piz
yY5VgHCsflVXLCgYIrY3WUhhnFNhHcNJ1hlEfWdfTPNcoDPmsqxjILLSvGJt3NElD6fMglt8RqLC
1hXFmYnlIDBWqe33rKvmNc62uITA5gHPgyIaljHn0tD1weM2pJdjWKZxk3IShcDMM+agUatoQfb7
opYBS95dYLT32Ry0M6PDzpcIVs0OIITB8YbcmySv1eJQaBPVqcObtjOtDrAb0zjT5eX0y2PvhIkZ
KOyMTBEJ/tsf52gOx7Gh0nhCYEjpKwWsR4bUJ0ciTjnMaH1ho74oBMw+Av5ch65yGRU7EJ8pBeP/
UULVbC6JQn34uco7OfU3flcWtkP8i9uToyiebT0w09iT7OUk2k5yqnLNh3EPFbpTJ3IF+GBtFTgV
hWmamyd1N6WV8eYt3/bQZhcZxuRj937OSIbUPrd/F6zyiFseCk7lI7tEr0H6rzPiAYoH+puWiuBa
awQf569JjzQJHSfhWRbrWcqXFNw2qUM4VdgAdcND0wsatCjYLY/50BbLxi9H6NsSvsKs6kIll6RA
lavmYYaBQB6AamlM28x95okNXrV8X8laxqkJRc1GIpLqIpS8S/Zx5iujYD1uRAnXCwOac78Sfet2
095JcuFZ2Sm3sMVUfzJ5EGDedi/Cx56I1DmVPkNwsp4wxvaNoMkQA6z3EbLEdokaEG8wyrxlvKR1
pArUbjRkPaWz6xtZuVNEO6EQeJEwo4sU8aUVzmXAxn5vFkd0JkLgmAdfJq/2IRz4aHBo9XpZIgsP
VPwVn3vPWPaoZ1njAee+Q5/6OWgxx9sz0k9NGgZX6+GNpRBLeguZhOkx7lMJR3ZIiy1YjQ625IOr
snH06jxfL6hNV0s2BIpwGAs3ek2sVGCHX0erNok9fbNg9dE6chh2xuKe/qBuzlKbLP1cNXj/7Hy+
oQ6kGE/tfMpNbaCNWjw6YRUKwHDCmB7I7SG6VlCATLVkve8QgkJl83RWLErqVs/P+rsiAiyd8Qg+
L8KD54xiQhqBtB2bslqBbj4BYRRXTkwnUd0LbwXARFEOt6T2+sCPAxv+PiSz7CFLsCLPtAs5xatF
O8W/Zcg/eIuL9Zz7Nx87TSe+Ao7iRUzYpOxfosCMA8UFSY1l3/W4ATm/ToBxUIrXJq4LXmU8W1cb
7kpmuQ/KZhOPs4is2wei+0hHlPRF3ZDDcHS9b89M9nyFY/+BhpoMKPrtis6wA4Q63HA0WGVCI5ms
hJymgwm3VAS9BYnuOZFB9gRn/48NlLXaAK028vS5W8NF+h8TYePKCr16KQBFRmSmUipg/ji/0JxW
LjX3up3VcvS6W4WD1wrKQ86jnuD4mAzETNIdV/eu5DYDiTcvrUzcxQbKC9lz53l+TGstzIY+Ycdf
3+VsRybYAGl0YXIX5i2/BXkwojLW4XRrT3aY3AC3cYHIkzsx+V8E9+Hn7xm4LcUWXfUiFOKBzT6l
mTuJmyrdldNqdqaW3xPMj3AO5GeBWZGPjOHMxlGXoOtUtTO/2xo1GX5qNuJ1iRhRwLPMnhVRO4H7
uyMnQJqIb683X4A3NVdHGHP8XH+bVnyeLcyujzJrEgRsu0iJvirU/aStkhdpiS6H532DQTrwzWLN
1lUPvRwuwoLboAIaT5bW3sdFBzBsTQhjk1Mhx2I5vPsnzegUXVhls6xq9dveSeB04hsqKykCWJ7V
WhAXVgCOCqObts+V/fHfT14/5AhrVOpHa77DVdbSqqK9wEOvL7R//HmsaXdKUEYHB5LTK/OtaNue
ZW8KhNlyNIisfQrtk7ZSFMiE03A35+MeaJlDyhq9E+t5efosX2fwntlsY4uRhtK3DI8KfH+Wmu2A
wNcMzG490rQxAWMpjGl/MjSc8BT53ZTUz4zlfNla9Iqi9PW/nuQOPJNN7l+LDYinO2iNUuYSvRVz
YJqTtZ7E1GLJ8WNhAdanKlOflk+X0GmAxRPLJ9/+xaI3LCMYsgv62GQhbNoNrvyidPOBDMIZ8bkb
KA9wsW4qOBOqS7zy+r2m967Mxd0S32Vj+hPSOm2ZOWEWtITr2dJKxTSmpvKWzjBejWDBVKknLYvO
3Ovlha2jHlu2ZMiVA7HDuH27h8AMkV9kjnwL+3WNSf7vwRXLq2E88Dg6u3q2byZlyUf3JJRRrrPS
Nizk9AFWCyTc7Hk4hpep8teNcHRYzAF4ecf4AYRgwo7OGnXi+VQ4w6ShRUxv6NfDH2MSlxNzLcFK
YCC2dvXKQ1jYu/A2CbrItSPZgXf+XzpFcXxe6rKVQSdGV/b1H+AfiANmMTOx8WEmwhraNcQwKUXK
qlVnBkolVFwPWT7iQAJsT9PSCWjxrtcVvRlZtTarWaOKjGpxvSs6pNAo/l8zOJhBujq8y0IjzcBb
GCo0YTfzQxalTSHBuRpLZqU50Njd2bQYynuOKFeFcFSg4nWuegVH2yHNT3ZoDYg9KfQGGpyOLRjr
CbACrZ9PLyrNz+eg+6ETWrCrgzsFChKi7EuIxGdkI829sKYGlczoN+pfEWaQub6lEUf/fv1DKG3V
agRiaO+EQhA2V11P2mjzpzrYH3MtVVLFPgkCxMrrNtqU59bEAZWKa+p4PWUmU+SgtnhrQP3LRosj
3c7+zhx0XyonNtlRyw/DzJXMOc+DOI4a0Q2OSpeYwY8pxdr4xG2Lfox7KlqcNjapR7rc3vYc2yJx
b+0Y2fFC4YsoGrPf1ihFB9j315kgMcy/PkVnZUTGXvAoePNnGkJX61LdkQWgE95egaLFdHpUmhgW
NXPOTvf2n2IdjsVaCxkAWRrKW96WdYdKQQPpugEtEoY3kRTOMD3DbK+lP1bEvW8H5eHPyUQVpS7j
S2SmIP6HMdKYjdBAgggvgDuzhX/cjLv6Li/TS7yGdq6LC/Blvb8NkoAu8cizbYg3CGRQ3aikjyRq
7sULRPYp55hIKXjRGdnXt51/gttWSWtRCDtx4R1KUo0+IiHyOX7Azbg0I/VCmt/6d2rAPL7IY7Rq
VOa8Vy1tbGrUNCYD49VF74l3dA8h4TguSRkzcmkjKEsmsNuO4U5A77l2ZTcxUgn1wcUiPlHbEVEu
b4qEa3fswMmAJV8Kl6Pcghuoho8PdpQwwoxQcCzLtxejkZgTHn2aZodnxo6A824ZuzfNZjhWz3Lo
CM8Y/P23sZDRPp0BNxzZDRvchhh/BIKi36fMgzgavNppitI6FZGnlOLIzmQPS4j7rNp8QOVJPlf4
JInfzNt55FgW63bfk5uqVXzDTj8ApmsWZ8Y+dZL3xE6fG977p/LbdnCkOr0JNzpDKsz22LX1KVc5
9Qiki6qHJBHYGT0DF4GuJDlOydMhxjlWmdrhO1yrOqkfKAgyyVdETq5p8xByY3O87Cv6sAY4knhv
ZQ0Y7tTLRrOk0L63hULI206gurniJIDxkxDny7yyYmxT6m+oMNBzrAJv7B7FlXrp7JjuAVLPU54Q
TZ0okLkY9w6iGEYMZQm0i6PNO9q8/30YDa7aAqLBGQZ3G4D47rPzKt7sne1QV4NVmcIIdbKU+APE
ObNXkSe+St83rmhvL7mKb5pJ5n0PoLhkqISDaOfCz2I4DRzRj7VuagMSmzdHZOv/L+x6cX0n4HZD
sAd7oK6ZrMOrYV63+RzUzp3+dV8gheuVHi6NkLQVhLzapLSiyz4gYOZSxe+cQjXxYT2XF1mTcfQF
JHkSKzO5LIy7eA3PI1doPdS9KDByOzsxSv9Pt5cKE4FZjZnn7SOKKxZgrWR2S2RCd5GLLYWvrOFI
VH/5cGRmb4KzjOB50Jt7E0+WQXRg8wo+cH+ddQC6B4WoJ0KWI4fSjJFVhZZlNllC/qJJIQrpISpB
70bshYdNUB8iwjqTutQlVnq7nv3kTFWPpnTxihLm6wqiM2Y0Z9/mrINwFuQn/TAahs39/B4AK6vD
R8CDHwj8Rl6QA12zo39XFt380LkUJxTZD8AGNBxVJimN4m4qRby7LD2WiRp6bWhX7p7Oe6t3oUvX
uCAAc8WnFkfXXFDVQMdmGNO8juwuGYDw5LDqcW8iDhy3aoLdzCiGY7lNKWGePjvKttMaTL2qWTOK
Y36Lk8zOTgsPfSBrtshtE8OZ4cOMD8YQ1hbiFiYe1piT755CdZxrU4UbSABXAbCp42wAw1wVJohh
YxjeSOphFBzFiu9ZnD1O3HX6+hKj5bMSSDPjgDZakwl5qHpeghFt+yVS6Sg4UIsLUtrCJ9ECM/wX
8mMn0T41yFhdOxVacHtLq/tf0r0pIaraBNt3KL5PcjpIyVw6fXn/qZ28YIWqNG1lMMLgQeGF9U6Z
54u84E+8wAhtrp9j5sTbyAijCBVLvBtlHJNQuVORAmeV3xTdZpich1i7BiVyRNcjE82SgZ7XamAp
bNO1bP1/2Fmjxq04vDeA1tOWnNTvKnFc2tmnEJ8NeG0KRU4hYYCFtzyDnSXB7IXyQQuMJ0xTxMCq
SxjzjUlKH+gpVy+cnhVbRRdJl2OJS0lADAuJfeRV0eQLpLA9USY1wBxCYXtkjhvIE6hlFB1A+p5K
X/pRCPtTHZVm4L+gg05v4QuLhb+/T+2Fnglew5A62oVNaxfr1R3rqNIubbwBoEc/Gw2xfejbRbpM
pPt8xy2tgEFeqsVSsj3hvlqHmu3cZ6xdWm8ik2tCiOf8Tm9xiqK+gql+BJJfbdHZoxlvCG/0O+TA
6EMPyIV9NRqMZ+Pg1ZvD+1+t7niAUMu6FINczPkrNnHz6N5rd2NNkPpz5HTWCBoZNU44EI3ckW/4
tuN+2/xD1MYx9CWfAWJ2eHKPkyAPYMmj12cp2EcRicHS4jNQ0ywAkp2Os5BWoxPWyxB+DxbE2+6h
oJ5fazxfJ/0l/Y4EwEs4h8CxxftyPlfpejGQQ6j7GVB8h5fWOOs3mrBfk2p0lA9UMAjxDJVqVpID
9XQxLSUcfm/0Iptm0675XopH0EYVE4y7Xep+CP9/u8FKCbrhD8WJrIEjmufjiGI+mS5Nsg1mo2mR
SYJCRv2bniwM8KGX6GiUI72vJh55pyK0EdFtasSF7fpDuJmkJSctigRdDXi6FmT3dk/RmXw4E7cS
tYNJOrYfXlMVSFMxyLWyJjwsX0F/lqI8Yp+ykFhng6X/CfJxcFbbSiD0wU1CDrD29eJ3m4e/uV8P
4LejK8WJRpW/i+RavmeCU4N4rdFgzQWgSzktQdiOzwI5di/hqjiEJrfYtReH1g2vplM/WHNENcN/
i7GW7iWtgwE4Ae6mS6Dtn1EsXlUUJhkzn+WVUxjPxSlUZBrMVXqFGFEl0qLThBZUREo8hf1fnVuX
1CZnWGYITAvI7DzjxEQ5Gvf6h1OCfoahY+hyPxYgOzQWpfQXpiuAMFP5CAQgAnLIYo9k+ftdMR6M
wZdfbRGtmDhm74x5SC7835Yq8eKceNiTVS8w61h0wH0X9zxotweavnpQseEQH2rxFN6MWd4V5TLI
IH9NSCE8uzyDxJU9npSRJj4OkrxQLF3k0jcOqfJUsDs9tbTLgALzQjnfOKispNTnyw8Aov8x+BEJ
I7r/1RUrcrgeJ48vQ7F1R+FvM2PAYkcjF+x8RCjR2fLlSgGPIvAKp5LBFiZHCiTe7DNiCvaJiQRg
aKNLn7Y1S+1xJApSCTYiHVYqAam4MVZr0LV1hL/EZK2DI0rvhJEMIb42uNK/hdL0bqrGSI4jbUQQ
dNMGMwXoto9cOLMc8H7FJRnk5UYMohO5A798hFs5f3unufB8LJtSRUmSGoL5c/RTda4IeHXo95Qh
HXs7fWcwqlbNCG2JiCvVZ/UB/PX2HwQC9yVpCUIQOZlG31noOn9diTg5XsEkD2FgW8PNoTz0pImL
it6UUacxoFQNDVY6SQLSbpf23HHFi6soMRyqBrZixvLN1aTOVYcXLyPxTCMo7XZB+8hi8et2+NdS
NBDkMuz+fgM7cy8s019PICzEqwkIYV14CsHBYJWW+hrlTAg9k1aTPAax3Rt5g76zFolmYi0bvAOb
D6Wj+bbha1vZTR/jXeabQh+62bnsc+IC5my4xYNnEmDh/u56ZzwUVv5dC9OXPE+2OBupbtH2WZHa
mncMByRhrrjVTOkSVG22urFTLwTvlLPojjYlHIKUKRWsW/oU9BjApUoM9TvBxha1MuvnopU+VETP
eAD46IR8EsSR0HZ3fPFsuV1/VnOhoBnWcM8aOu9cZ1jHfkkzs8O6TgWr2EtuMID+PwB0OYE3SKOP
DLv0rLDfqlZ+LZw0ntZn0VXZ6hm2G1kOE5XKwTUxyqA3AQkPZWuD/SWAqq/f4t4R05TThedqRstz
93yBIY0N1VejSBkzuXbx8UgLUbciyIJrChuvh6qMw4A8HrE6dOF634SaI7NXCU3bZ0YKUQbpSvyk
nmrbAbWpJEYjk/T2VO31eY6x/RtRRHnQ5qKwiWOi1hZP2nZrbtbIm3GYx83KSHa/e8ZB8XekmSyK
J7ICceXWPlsFnQDBVeMJjZ7bTE6//AbzCMxmJ2b6lZ/Xd55aqUihUR+2o35h66Ac4hIG9sJChz9X
SIkueuQoF69nEOR7hGAVmsgvLSahaY7nd4AfgrXfp6Vo2ZXd/Fxw2BmQSwryO59pVCse6HI2myh8
u7SLhWBHAQ400G/gEIv/9MBkUR8K2s828fbK2/sIZRmhasJPhJ8bV3t4WMcBPtw1bGr0VORdD3Ae
zBqrOf57a21duMsu29Vd9k0p9SMN4kcSQ7QSWomf1eIR2MTo3neYvU7tO0iBmCTrq3jeoB/ktAIR
HZ7Vf9EqWvX6qdD689S8YwEOKXYFPkAiyRwCZVbHq3yb5PT1gCFQyvn2oaVnG3PKHgBTIuwWUQya
Z8NO4GbPvQWQ479n0msiCP95/e6QwvGQRH2ZxRxnOCrra2T0GoQ+XVUBTPcZV+grXa8RgOn4MOwD
2VCQ8yv/P0Z1YDjkRalH2G6rxKQMO0Ii5i54C/hx4zpqfnDxtFF1tOZZfpTMK80f34NClSEtNpLt
BziW80Mo+2ExgFjWpNJU1+c4A8A4IwFsLEEbbrIBKZ+0Mxd4cc6I2bpoIdJSK55vThHD85aE1Tfe
7KnVc614PrweOKdN1MYXNXpd+HCE8awUUEgBCNKmmruO4WGgTSqrti7K5h1CWOMCnv/2bdXR+Vp8
LR9HjODUpWK3B81D2QAPDdi4bZ3zas+UXi1AdjQVnB1oHIxHJuiwF2Nc0qfhUiqZPHcjEHuJbva5
Zm/86YvprT6+R9eLV3CZksoYzdykQnQ4aPCpsom5K5l0Wsro330IODbeJTgFoaUq6MrN1ekIbdRG
ifhyEEt8pr8lRpA1NtZpYkA5bd0wCs13hjzOsB2thaBHnkoXkl3n3gs+a++ogiOWEE5UJ5CNVduz
1vgz/tT+I/OS/5Kl+KvOYmxGE5d6I7pjSi+pRwA41Oufxgruw5RM2Mb01E0oUdHKiXr65VP2IHLG
YUXJxWS74bA2OOksgGPrUjMJGAcIfG82vhYRar9AKP4+Ilo0pqtbbZ/FPG4T+9Yv7yi6GALm1euP
xETHlz/C+kJ7WlORvZtjfV3BysnACBcetEqHOA1u+on5BDpeSAmgTwuD7EOgQ8nZyoKITkuHIYDG
oeOldLOJfck+Bq4oCjro98wiEpv9zWKuORvphpnoazPvsOERgx2ovPwfVUPac3N6APixqdq6xOMY
z10h6kg3fdiraHdm0GV/SdDkvmXjVZPXZ+4jy6FFw74dTcIwGs7XsrFMq0ZKEK/5TeQD0YGwcaF1
kSmMwn9UmKH2qzKbGkg81UlrZk51pzXfu2HP3QfLsAh+UtNDMSoXAaeauNwjRxbzCMVqE0sKKNXe
B9xs+pSMR8zd7mZ+8LBL6Nugb9sJOMTrFeTVY7E00B+ApVzbv0yBa+a0VIwG0aoo0ISMRmrol2Uu
JyDD2qB+hJNG0TR4TDCVUowBUxJ/OEFXdrY+5rH7EUfOFuRzNz+M5K5xvzLLkcEO9+sNyiXvIwaD
xXV9SeLAg8V9yC2e18TE2eK7eMqHLEcBR7OuADn5TY73VZ8R0adGEAGKvS7aLUQqaiyhMCN+xkyK
1UBnpRiKxdXoiEt1SfhX27Fs4y8gNEFd0FDKdlIiI2I9QqurKkGz3HivRmml0xaU3tnGUMCpR+Bk
h75w47H5U7ON3/2P3y2gg4VTaf5aZNt3Z+PMs9fbDW+TXEwtenQvCo+Y1x2tz3ScZ33mzGaMJ22e
ghUu97Pwfd3cV3oNdEZ2daWq1Ytj+LqCdJzYazvdAFpcBe7WJzOsN49oJedfLg7/cn9uOFlonT1/
UpCg2Ahv06Y1UbuZX/Z3SEswTeixI9SVUm7KXvfkenHLGxnNNNHSsjCDXnMW4XIIQwUWB3R+KL01
SVy/UAAUSzYFWpYTp8xYoCzPDsSVfcWwhs8LDgyu0PSltIv20Mt9crAHGq9+H0cLz847gONEGSo6
Ip1qJnuD2m7r3woumTHlYxom7wDlt2MLi/2f3qnTrhRwvzxmspG+BmFM+m8kPzmHehTk2WVejLHe
1MK2zlfgpIOPbYXpMmWcgxjG1WJyU4W17jMr+htDfMXjNK3DYfMTnobIjxdwLauwjO76SVKU86B/
o8f/bb1IA2vD2oEwdPsXC7f6/CLTd5Z4yMU0VSPSBtWSAmH2GcJPyV2oLd/T/TuUvXqEKzHG2NXU
aYMDF0KYcQVdIUdF8mtvwk6AjG4365DlJxJgaLHUf1JTsXb0LOjhM7ZQdGCv5gijpZNIUJxGtF5Z
Im2IkwmbEwcZFemDKguganQo/TULy43peAca5uGxw8wQQMYZlnIUuFoo02S1AKN3UigrJM/FoMJP
Ss7wYfjpvOlQaTKjfJ8HKrfDeufSrv4cMeGhrufFP00hkp+CTBra3pQnu12fEgwY5jzK4l+a8sJS
vl0rDwOs6cNygaRbHtHRMyk7zsTD1/KbUymZkETDBMuDAUVZiP3Chql19FADGPD5AGMrLndHExc+
s7X60HxSKIvP4brQLyvl0VinB1BiimUs3IF8J8Q+CGb8FKDXs+APrFe/KVku75PeMTbRwjirAjMa
K/g4DF4NGsxlMWnd+5haWGSUR4p4daPKVpPTx9SmbC9DBiMm9dL3kIrVJ7NwfObwCK4igiJVr7HL
NRiAg2bbLvadah0QwTGQT6jIcbBFUdaHrfhPqMe0fdZ988F0Bz2QK9fT9BZtLW/LlJr5a4nUfn2z
WBsCbMcZMKNHL6GHz1oOvRw3PcWdmyFxW2jOiQT9woEkfrh8H/3e5iM4FJOx4XMCi+A9d2ZQ97KM
ixi8y4yff+U37bPXAvbK9+37F+J2Idl4glRizFjyx8areIjs5tZggnEdzgimcE6SLNL/VLMJTGcn
xJJdO+Vo+FilHOGGsX4qHcRwu9/IfWlOgSSdmhrmy2c4lBIhge7evyxDhsfhYBNcWipLxbf/WowF
xYXuF0nSKzNnEFD95sqBH8tn1KqdvlXW2Gukwr4h8gaWR+W1UBxfQIFtL2BNhcDZWG+7Ap2a4l2j
G2QAZWynMKpM9mvUTG1hs0uDe2evRrqdBK8QCWTnu/ORcL5DI61Qawj9DYTxBsgIMPIoiBidStp4
wjeaag/MrLzvnQOctr+Ipv28jGEUk2ORFUIBDRfAvYXH8DECTjYwCijK+4gXdyMYXTrXU8HfizVf
tUndfwtZRpCHfnYKj4s3Ku8GMpUX0Hd5Wv4A/1h6vyV1x6Sh6zvh81Mc5h0Lh0zi09QgISjNpxWJ
xx/KjDucbHjhsPQrYgrl8Im+OkaMnLhBJwz9oQFMom8ONhzf9cH2fMZbolDFeBu6WEvC9naWRMj1
ehWKjI61AdjGuKWl3dYxTnISwLQNd7h4DAfksK7Wt6eoCOh0j0SPf71RNb9nmsYx9XUY8vgImjmV
3BGG4DdLiKilkDBC0SJaEojrhmHyy78tpGOl9Czo5Z7M2fb/wtxmp0luh7OvhY4bs53VA7M9vFMR
sBAvZtMndm2HA2xKK/O6LcBadIxAy7HXjjv7Cl+3ArD+v67CueLALHSuh4ItEY4oDgjCRTS+8D5q
CJmMUvp9bv6VUDJRDA/EUwaY/FVtyv1/MQhY7zcbihn4yR02+nTpdVkHMiC0G0cV18/G6au7ZiRC
kv6CUIfuczYuv5qnlESgZlUSn8fk/1XrgSj4u924lx9DvxX/KK2jL4OrEe9tzp4F+XjTL3pKYLWM
n6elADur3vcWPE54PJJR976T6K4bY1sT4oxYWGzJ0cBk8q7vD5GxaWyidthkkARlzX99uBw7fbte
2uai12KgyPwjojbRMRZ0IPlU9nsWXvIL8o/LmfSnA0lO6TnBOCA1LvS3FDL846NS9FvA4++iucQz
lZGCAVdqkFdpBMPadFNK3ttbCx2AHvjKPZM+3vC2hYRRaWTubk8MG3GGeeHd+5cceKUtwuPyLdr6
jHcWnNKFpkVaUzQ7YlbvYE1an9klswnPTVdF9GwJi6lbBD/S6qHVkSY59UWNbF/cwJWaEzKV+JV6
5IXN7J1kvmvJLQBgtIItRRYC8qk1xb6cIpAq531HK1gvfnLQ0PJgLl5DiXWauwqzaGHDBD+5wbve
lYnRDuKjpfzDyeMWGhXprmjdro7LUK89qwWbH3MGui/2VZlFr9HNWIGs6alUc1bVKmJ+NEb7W2ul
DOpmbMBQZbloXj8hBkoHvYkqNFQhC2zo8Wv8TItQ3PGiJyzrzLIPzp6P092qcsze5ILBFPAyQYme
PNSExu4I7h6vKeo7eqIYLk0wZsFoFKBrXIC0LeumgXwMu4ATpFLjtWbXf/Q/SVVC9ivdMTensHqR
K2rYGPpodCGk4pkZVpz5cU6Ld9LcKNvHK1CbT5PM5207ZtokQqkPI1CVslmX6YRL2yCEDF24j/c7
8D8pOQt+Ug/IViAd6He0L29FLg6rqNlG5kfkBLQeuXxZNr+wFhGT5Y9ZPq8tnnDY3S6jtQfbgyFf
ztFgHmI3JHEIfdFBNh2ZFSD2h8oQ0N/SKQu6UlRAwz569OUDbft4rIOVDmnO+jpiuqq4yv/4LLfw
YF7mWgzoVw1ASAXptROjMVfeEXDNPxJRz1sL6ry0HKAkY2gkhxmQQMjzRJzG6iq9JK4A9K4cxLcm
e1m8yYNqp9GYFXQ3buFGjwmtHphqn1Q6GSNT4KFae0/x87Ayp3Zx7GVhSUsFPNWWVx8AdK9SA4A6
uCms+7/gET98kwTjAsd6U9CK1tvQ82GvngnDwCeywrKPxttSEhW6OnUjgXz5GXzh+AO6dNZzFc/E
NrjhQlFIqWfIWUVYFibQg2pnIICZxIbxtE/J2KmfWNT4mBX0eyslmKx+e/4+SWPsLHZ+fGWTZXaw
EgU7TuSI+0qWuids02kYAeeq5PiG96HfhG+1nrAqapl7lTZLNT6dtv6nrnLXfVdd4s/Ut2QHM1Og
DkGlEsbpW7TdJl6poWDdt91b9F694gkGzmtdShjddvWAcDyVjyulETHBFI4h7edFPg7YEql9MMXy
P/sLP/wMzV/ewbGOtcr4z/l0EFTsvspI+STvgmE+frD3vqDWhtpCn73yqu/unU3BiZSGT+vGbJyy
sIzyrlK5N93F63tOgpYM9/Hcl2LYTF9GHFF89A/13QRj6mOvfP5WpozQhax7KTIaEuGWx7TKxbyC
vVelMck/X5/zpMJasr8YNEfOO2kyYOHs4Dbr9WxCbwzvf+qxZK1vaxXWvbc5rB4qOv1eRg7G4aCF
SVwzRqYX3O50k6uJ9i2nXEm/0GMYPgDwx7O4pJGdkWStwegDWfpaHf0wTuPEB9Gmxsv4SkGJ3hKy
LRdy4GtNaNq/pJIddwILWhYeBnNegd/tOF+FWPeBIAJ2KQY24N1SrF5ZXVoJMzO+8t35RzrcGGUw
Gtq1FG/J6eIVKroy84rTQD2NX6p3OUxK+lPDGsSeOQuE8vS5L7QWwblyChHTTZmo7MMslfUCL8YD
WttzOXOP4sIuvNvd7GyGCkKv6bkr5nqL7eCPF9DFdFpVuIJLPfiaWr5flIah+92uq8KSC3bfd4SH
LCtjfw7CYCnCQaHKw+HtWGZ0c6GYaQOD/8cqYVNkrKnIHzNlV/XHnPL+YYq0JO+vLJPHZmNCeGeR
QlkGiI8BbnlwJSs0mMAjgyP7hlsHLhFmM1v2ZttTnqnjQ+494aiAi+TkCAwvFk+/rHYaRw1SMbxT
ZAcjXmVm1TWiT8nYf/Rqq8vPu+lFj10y4TU214q1eHzWBQ8GtZLPouanyxQq3IGlBmIB8k1BikWN
9m7TdCeioh714dkMcXupxLHg4V21U400b78DwRMfONvnohb7cWgDY8m1q2S/eeDv5VPLRGxw+ys6
bca42A3t071qyz68Jg48qv2sEkvfHYQOkhG76ePGFV5BgfC4phMBU9vBYk+rd34S1psnUouMycUB
0SnGsEQNwpSECPnVWmTvbhm50UArqVv6BtgYYH7GlYBgIza0gY4K3EHRAohbGZFzt0Xyy12c9rFb
3w66pr9feeqWsWXn/AnnABeKWB4FLZY7K78JCuoCpmPE3nejQTSIfdT8pPIOz/cKzRNbZzFgX1e9
zDITVGopkkbJk6XBLzlD+rxuHT6kHHrhNYBP0RhGj4hIFdKLvCcsxRrD6lWVpcVUktrNB7yq+ING
wR9loDsnxTthO3Z/2nPHqyM+P9x6qxOZ/lYq1E3poJ1wwKddQWucZYVIEBdTWDCwDUessWbju+km
1ackei8zAcsNlDaDGBnPMCiBJGNun8a0eWcyDXWdRjcLsoKVUnbRYBDhzhih6e/uQtldBmUfL5Pi
u/cg3qklBRAG9VAqeNEE9zgfZ+g3upTV5J0L/IaY2JC2wmwhGY8HZ4ssw26VgwbBEHx7UTOXwJ9X
wWo7bUZrncW5Daq3B5tX9Bro6sdSHfGpDwWw68I6E6jZTTsZundNab6kIlqk0lCbqAbOnIHueluc
bPOn0WWVTPlau34ghqB30lLsJuWnhXGifeQ3HLpCBm2nvE/jHp8aXuFxML+KY/RJ3o2sMFnL4Soq
zPQ7YGkPw3KLVV99IcZ6TUxV2wLktoRW75OY4oJStNtWzyFmGrFNlRRNBNHFbxEagzK8i7bK+GhB
MMZrlIXoaHD2egFyKt/SmHEEwo6yPyAELLPEi2wuQPGT/O9h0VLXrZkKDoMJv+ATK1SA9BmQkHrq
JaJZU3i5W8/DWSnqhKOb7kvSRBYuE0NXmKAHCnqYXZArudSXgDdEA9IKqibcfNnRZoeIwvtUSbUL
V5v7SVIMkNM3xrdvwcyZ0cct718trLJoCA9Ky8TaVjEk1EWSBpqGLY548X6q5Tpf/Q4iMooj1M0C
dgR/wWMz3EuNEDtxtCmhQnW2n1hQBSpL1MkaIRevBHdKkT5FAK7ZgZbXWItc1Dz+d0ZgsZ52uu10
ucMaKxFZwwGuj+fz7hJstIkCvDrEpt1VPfHRugrICi7sXw+WPVqCWBhwUIh8hP7/9Dix7+zizkFb
QYxu5bZjDJnilxaRk3GS5Qv570+AWi/1O9RuK32mpy8OLcFn4QNzc9nlFceaKOiHzhLUZsWTg0N5
7QszSAsZzo0gP+55qMUAXtR1cpNEIxZwD66+MyX6XcT/lat+MpyGQ/19cA5i6T4O+VRNx+EiQ8Sc
P0/6F5MKJkAcQ5S4JqWN+1bteNb+SwED+k7816JQ+0vT0EB259BmIaekh+Sl9ENpdJx1VStqHN34
XOHtQcxBVqUc9tCxSU/FHnkFAdu3h1XYlyjjXubcMdlsMTmnb0i48ejuIzKIfE3t49VRm6AUlZ+o
fTaVoRiteZcriG4nT5y4Kd3BUCtXCcFnCBRWBAYA1bAiQK+IO4uV++bNJqctsuIqtheaHY8W70/P
v1+KnXcv9/R/0yEbT2h8ZoUEciCsssvkJ78Ezq76lR6X8a7Z9DuCdKgycOMyVQt4NHDTCp3E6Pj2
3VE7vly62K8+6cKL+XwG/Wcml3Qi2x7NHZeY/y1iXNHUaM/nLi9FFc74Rf/OcZKUJhmPlFr78ILs
WyBwF79VWxrxU7wVW9YfwhVe/9BJjp+n56zRF+PEqx7G6MXQaI+6pCnDa/IXd1ngB+E68xFrPklw
pueXGHHiZft4MkKwUIm7QgZreBL2Ut68bqWW6tiXIOi49VOk4ie8/slOyrs72EnP1SBLfM17vCAr
AialJ9M2vbUysBEmZNbKoiJAv3eAPZAIlezPqZCRYVXoFzPt6UfD/T89NcFmJTQlmLZsMYR8USoo
km06Sr4LunwHiuNKA5f8OKyC4TaKLgfCPU0KSzhqN0030Ci1TYt5UpPM6kAqry6uIXPrcVOVODpU
GNrxt/Gv4i5L9c++cTuUA5k0t3+pn8j/uIw72MLWVlla/1tQ83aRGD7jkpV3ELCO1g+os6JZAdg2
ONr7k9aZFa4nLw9VPy1MdX8JSb5TpCIwvuNE7/ccgIH2OYM7a7Tg43GuOGTiKUNNHdQ6x2senZmu
MHXVrqjYdYq4alt4PXZwpo/KWMkHEXAH6qqJuKI6CtPLYYSjw+QSLhVpNwpmj67C6m/Ihgc8bZV6
fJaEfGcz+FF/oPE+NKSaZXuHpQ6VkCJ7XcKgmr8qq3Zt8jJ8UqyqKC9j+CKc5724Y3jOKttBPBhO
klb+wELrJqSMmQOR0aJfrvIkT7Y0/dLRTzFX9rkOqtITlnyEpQTSoFq6LkxQNNFEh7ZdgYZE/Kjp
xz1UuJ8/4GEPLfIhpqQ9+Us9sHKIg1QL/U3FdGi+OA3Nxrc7s08gRU3qaeMkDEFzwAW6elQ2YvUi
TRUcwqH+3sFFoFogGHif6p/oPDcyPwXjKLRwBspVjgvu5okPzEENFtS9U9bkHFFcUwJhX/6zQ0jj
FdUdAvI+QFsMZGN7LK8a2VP/XRGRNuAhDadVqKICzSLsW2RSFa9kTE8aJW5loljhatVJ3gr2cssv
rF4OV+Q1ybfBiGWNvBQ8AvlqUUxn7aDRVHtFd0sDCpJw82WjDfflvH9G7T2NrwezqSwxyQwscmBI
GG4sHxQxIzyow14CIDaeJUy9XpGgRqRMMMw4FVOS73P6oB+bsKqMa5lrmh/2O1R8UnIIMqluOPxN
C/eTdq1xK3rNTZQ18zvuuUQXBg6Xahrm9qPpzn1XEEIXo1vYYq2y0nNgWi8ApSlcUJiZntyevgKK
hCceIuxlsvDy6kg2yFsZCnCfV0eHaMpDmjLr6NT0kSmSQ9HRgC5orfQSc7pRLHFMxcp11VY+f6ts
C+jFF1ZeClPHjKLUyzUuTFkhiZph+sgygXiy9Kiiq11qECWSR1m6BAgtjJ0HPgdz0ObACxPTfD7b
uPZ97kQKreWhLi2+s1mCcCHIiOUsxxxeeQgnMSMN2JBdlzMiEW9rdeQXvoa+sP1EJzROugr0fnEI
1dtWpjsKA6vzcQo+ZAviTNBthwSuqHDGjsBBzcGZh0QW8JLiollVo9Bwbu0NUqyQTdComnkFkpYz
duklGuKd2gD4q/10fRGGnaP8SFebWnLLXaoZyCLqf5a4sF6jXWbFASJtObUuzlsGFh9wL/QsSpou
7oayB68WpyIRvWThKjaxtPNzfL3phpEkkviKJfwmOZTG9aiL+Iz//KsD0UkpMlbVxSyYRRpy5v+k
Nj/rRxm1PsYrOhKZ/gAvvR7sCACNcNuTdDbWhohJJxDL6AggjqIWRLE3eQK2Lh0qfTiTeTVz5MSa
gCg+wwJ8FhHJPz/vwWfKMkFSHGT5OSbH5jZ6dSKOkjnRH80+5btW4pL7719tPGeaYgt6kI59+XbN
fPkkqRIrHvAxU3ff2/6SPCAZsp9v9zKmlf15kuZavqSLLNdkBLqe6q8ZsXfyHZMMng/KoiQI5WlD
LKdJpe9TP2zPt2Eo1VFiGCtY4PFke/bLEMjSCIgth9ooJweQFWvO+LKNH4K3YD+dC+HgZQUprUfE
2dFIYhT3bfxmnrqD8HThV1SGxHaqqI+/xKE/BRikHHumzOmasWpFC/u2I8QHikRXXtIFjrt/c7Jw
POlXbU+ogy81nPDcYgrBdXoixzjYP1+s8ODsUYBnrvNSxVsTqr/6she6zqrVwmH7VowGa4M9Z96p
JfW3CYo/QtVYJfAk7G4r1IKpDx7VfaVP2AMVn/h2gO3a5odZTeVL5/y3ay/teF8C/fRch5piMn+i
cENTIGirKJyLWKXuHkr0w2+h43PCb4sRy12gSH3DnPW47Xu3s6YX5r6oJaEHq4OmDLqmA+wFt3F/
O9l8aFijP+hUS4ErDRpwcDfEVYgwyj1YSJH2U47kaKn97fbKoSTUUOFHrLRhP3vVt9FsnZ1naIFU
cbbAep27hlYZIOjZuuN0xlUj2ewvy+0dgcP/WrwYn4rfdYzHpsYrvgn1Wzy6J2JzvWAUeYKftHKk
ukeqoPvn5tYhNjJ+Vt7Jkl4tQ32QjyhpNKP4j/GNKdOeoY37z57qr28byjHpfGtSPsDNjwsBOpqG
tBc4h4mhAtUvCMZMKE7vwLCTl47Sxn4Jf53XPpFd0IZUt23kecHibTKGE3fCI3l6CLtkahqKXsko
D1sqeRfshA5ER6Fa1TLo5/Aqzq5jF9e2Q6f1V5cC4GFepGvDzrX63/QRT0c2HqXCGdURDbq9u2o1
R5coclFo4Er0V3RkaJ3ooRUpAT3ofZjs02/DzG6SoQrjzuLd0LF4aLREoRtKIoARSkLX8rCkrjnI
AGqpXneP2nns5xjQJjtx8/2Jm/RQ2uKFv0is5b14dm5OFy53M1ZMGk09Xb83TYAH29JsThMpkjQu
STuEEeofiF+TOkJi9MOcFwDbanUQ2GROLW/+Ej9qHuTCjmrBd5X1njX0CpogW1AaSD4hKyzIZ1eB
71GR/14e3m6nZlzCwgBhq9EvxlgOCN+xxyW9qlrQPeNn0f5W/vHwyELGH0HR9UxwTk+KdLM++8qG
6MYsUTZ7reOSipKisp3MyzqIK4f0NbWhTZ98RbGWImLwOetUtGzrKuuzklyeiKflSmwVxsvcdQeM
VYJ+jMFiI3ZVe9zqGxj6dexu6Sc9F0M1IUvsqMvICfjGQcneU6I4IeIYYwlmCpWiyKssq9Kzn/dq
cX9jMYmyEGzPxKiVkvWVP4VbvKzCE4xTXJcGN0WPUT5putC6C1ITYPyZU++e2hEQUO369XeRbuDQ
c+m4qmee9bayAXsvdlSTUQOjWZGsf9kUVrqmbttcPlSIiI4PPHAmaCO7OZcRQEAR/zG3SGD/1Unz
QCm9btLy3zUPojLwKiH4gLPgFjX79mIkcJIiGCnwCE9pgChu8k5iViaPs4gQtklcLk2vAroKBkFu
sEOP5x4NWFGUAOBHHQknxmhek+NY+cnfKmmdf0Wosx6M0wYkoxi0lAvkhDH6ggakH4sYKB+XirUN
Mo7kR0MQ9tLgAlyyf6CnKIPVVATIX53IIu1fKLIGCiYRj2MNUR9sN5tPp5WdjtZ8CjhE1CmZGqmN
9Yt6KlgoMkZPmXGgSiKYlQ2Z9OpefQTz7E1kRTT4DVPobvzpqbcWZvcF8keWAHQyynF2kNpk/0w/
FUYs6h7nUyogUmDtpKmKCvQENZn+x5deHxI2rZoDa30r0Q2V5Ka5Fz3/BUwuCvQY+iuJuSBSBGBl
UKpHCAa5LfAnLR7E5UTSyW5pr/TQEMZbtyHamS1/ECqHzxoJXpo0/B+qi2Y4SmjOcfxnfVuppfK8
Ah51LdB5DRP27BsZVYeHUvhk7DbKV5GandtpFd/KZNZ2gDXzuAMC6WgQbhdZZwupiQAvq/S2k8IX
ua5DtcK23lQuqVtjVPke9kS1zXESUbR4aTriGLXqy/guYG9felYHOIaKfoG2p6ChYEYEjt2+vSRm
j+VYOTwZHUKprAn8rHJODxrmnIvv9kHaPqXDDUKMGZCTOPU5iuQ7iNRNFgRWc5fhW2OyoEPmN8zf
9InzMtlC0HYaCP2KDOtvppgZfapSn4qJnfJnzmAe8pQ4S8DQ2OxV0xyps23dvuyxdXjlRfPLiRl3
norhPPxnWYsIG9Oya9LEWK/+SmIf1cJLEPD/ysHXXTK1nsNaV5yVU9LwfjlaHT/6BewYw4CO6eHY
7F2KWBsD6IxPCHIHPQtwxU2IcTMLyqYHIiODeUYgQdQxxj4mdNDAHHd367oFHfort4M4DcYEeCe/
9yabcjQTCv0hg2BlJ/6VFrX8lDHRXgIBR7Q0Nuw80c0xUk3giftuvq4DREWJWqG4VM287792RLEM
tO/XqtV3p6xGcxVIkatPdvT2k7yEEDg6tyhCCpYkg+DlkdhGGyCeVwitEcMTrkYEfSTNj1bFYIYa
F0TIUAZ6cdh4Yipdc4lJGilloZ+98Qz2apWRC4k6+AX728Wl10wDZQm1XWANJLQrdk5l83mHvZGO
rUbLHwkQq1ECBSOBsWOpIYaUCKqKAy+W1smvDY497bMCko5g2s/DbjXXJnal1Qj5rx9aq1Za9FKd
nYNYDcC4tl/jF6xhguLjCx/JaWhTIiUmZ3kAYQquhm4MA3RVKtwTdpS+BvQi0rCJU0SYnAMIA9EB
zrQsRnb0NMsoHrVlWdL+mqKY8XBlTvDMBeaDqomfLUdBNsioceqltKLIQOc0zYYsQfBH2r0KKG0z
EmKPzxjWq7U2lIzdPWfNLpzKoIri23JGfGtwFh7q4cjc3A0A4YTxWDnouVRHRdgrZDCZnKfdRfcG
P7CX74rZkIJq9deXRNB1YrRYkLJLKDcIY5FCebUJdAdA9sARTvTqZqN6Lf07mmMOZF5WgFgB4R/S
nGOCBgdGXPUtinVs6LPVTniPrqGPInwCNheJG77p30t1HvM3SSbgZruEZk8dnD8CdSl5iD6YMa/J
D9OXBcg/Gms/hhhJlODWpf7PWcbDFutBuWIxFQjfBuFMcMfYUgkW8Hz+rSAeig9EKxohN7plfzDx
c3OEgtfIoU3zG9obKaL1BfH/FWJT+CfqCEItsyQ+1pntFAyyIkTlss4pOFxB6LPq+h79LjJP6XKC
cw3MMeh/hGAeo5yo23iItyyrUzvRB8qY98GToydw3aB51XluPFARf4ddjnzENEcKfZUFvh2wDuZj
KFlM3EnQ4rIa8GmCEEAoHZ7MAhKnfx+La0BnhErrsWXmuYqOc1QtZFWIAQMFoeO/KXYePMpQHodR
IjIPRDOa/1rt+FLfK5PqFeIYTaDweaxg/ZA2LDp8d4hbNeJlsBM7Z39ZXBQp7YZyU+rGlNWzJ8k1
Z7ACX1FdZ6C12UI1jTGZH4vPl28YFjGzJaoQVgyCSp5pw4Z7hmRV+uszfvcBxCkxvouv1mIcZ96f
8UrvWMBc3ArSt8XvvtM7FaNrv9FgzPhXT9i0YkowaOX43+HU/Dv2u7ezsFmqhjPfWGEqIVne7Z3B
bgf6Vf0lW7jvAXWG2lO40JVmLA3Xwy4mzMye98oWH+sosz8KuXR6Yhwlw+Sj/1qm1mEdLP+BNcj6
2kU9akkVvMi7M7tuY0RLuXRffdOFYutqFRJYiLO3KNTBe9v6o+Um2Dq7oqNTX6hopgiJNnVsXL8D
WhVMWiCcwgNYeAYgXXZSIrYejP+vlhPCeWVAlM96WhWPmnQz5Q/yOlybUQlO8E5zYfRqfyuRleCo
8uQ1UH8q+g172f1fAmqF6sUzxe646Jz+Ivm5GmR6g1jqDdOsE8w+S+2mPYKr38wAteBanDY6ml/U
QXDRIwibmv7UHkI8Ag0gipgdJnDLkIz+mY4cBONGLK0KW6l5XJZtZkZmJP3FSM1w6ZC2/98NW3+I
xJ957nO5hdd2osVADowtogVOvm/U7GvSBmhoLd77e9QjUJvehXT2mk0c6YVLwUbBsDtYxNvTo2UM
c4dPRgkTkiJxFlp+CXg6H2G1aX80dGL9pFUiU210x0n/AaZ/A4ff2c2RdwvZ9CRHWLv68Rm2W+li
CS4a7roSwTEERxOaAOWDMX3KZmjS6LtbypZjAlz1yo3fQJO3kc4jRdLgjXGN+HaF39ZjFQ8H1mMo
TNrrSaujRMW7qtAg9T5m9Pz5oyvYY8UXmc0KjCFWkX12SJICbAM9/OgSkE01+9vTg8mRvpFZE4vU
ZzyljNk1P0dpcuokkjNoY/UyDaUffiufWgpeSaqxxUN1kotJkx34W5l73AhGGqq2/XaKm6X038nJ
1P83XJgFvWAQ7vpQSq6dBnf0irL7kqIB/Ow9MwL1WLZTUVlTb09RuOEJ+qCniT8vmRcoQoLX5e/Z
WAiAXV2avhfN9IUv2TKyj83437iZVMY4n20xZmzm6pqAecoDrxoGBRwhX/Eo/sSettvVSYotkfoz
AL7pUNUJBaPZBb3+WmvzZImX84m0y+d9y4dwki2NNxOptVpj1DX7v4Ih3+aLPqvLqdT8ciEJr2AB
SPd54D8y/YriAZcfG+/wUMFfq2rLoJx51iU0ckGdQZ4nRYP0at/6iQHNKAsuVNFGv3WIOA4bDrUY
Hqx9y4lBPb5BpUX2WbLKTjXiTbUctliXqQxO16mXtkZ1ndwpkJqAhXZ2/mo3fJaTxC99S4MDW5yJ
5RgyM2/8VNFHDLOS0LuSaDH/GjYavzWzgL+ovklSoa1WLo/cKxC/fwgWAnblGIZnuy3oQgmwlDfp
PMNfRHNnoYN3U9jF/t+RMXfOhp2V9f1+9HpKUnxBJXNw2rp/VORLY0DRIzvvkxkgnhA4kXUqjExl
ETwqMuGdExDPpi1toobdFzW2D+IdgJM6ZBXwLG5sIOTjNK9oJP3Orq/NUQo8StZ8A8CaFE3Iqgi9
OeuIEx4sqHRH/xmfu6AepfpOPREv6ilv3OuGYu7PvBLBSJmkZiVPeAoyoGhgFza2pZlhE2fgzcn+
ZE+hqlbFYCL7RZG+bko+ksgYHCuae7MvNAOFYk/5cGpWqaujBIbAJ+XYo2e0c60XPRUY7TgnT+xa
NJKQZslxlzvpZqB2eiHlAh66xOcz2jqrxTRPe7eCqyQDVMSbLmGeNYudKx9Ja4h2mpUzlmn8lavK
Ed7WPZJQWIbczENuwjeyWJIGQqaFgTHCqXmNZhKPjBBnXlvKmcQQqTbp3KhCcZ7tqTkAo+mZisB2
2UMcyaVUyLyyKGBhAuZBbjxn4sO36Tnro9EXtiGP6wzKB94r7b2kdMQA29Y2TyH0x1iiAGLkdSO3
xPhS8xGTm3P0W6fc0ApO2NPvDdT9fXITJ9kUyNBJrKyCWAbM7dKGDLLq6qe9ItRqi82uhpUSqoM7
PU5fZk7AoJ9unKJlFD3WReSjYiw30JcVeJd+F0tdBUS+EX6KdGF+nzM1lKl74l58ODrtM62egzqF
LWFi9N2ZPyW8+7TPCSv+6tndQpQgtmPLCVEbkGaj7Scf8b7UrW87DHo0zj8QHJyYdWPaOTCHdS70
m7wbTkZA4C52K9EGOpeQBYyrYCCj963Ps2GPl9NSxOVh4nhsz+joNTihvCEungC4GYFgFDiowrEk
l4vkdq2T95oViUoygSit3wzDQszB0RJekU5mLIHBWa003yz9+un+FWGSsMm2uzHMVQZvkSkpGOvo
5pMybHEwgU5AjqIEKd+0jUe5FmEumnpkjqNybdBpj0a3O2pTK9rgfB8LWaIBqnJ6TfwcdEpSfmmm
ax6Vv0rl5smIcbUBIde2kZa+B19p69d4uuMmgrq1AIFp1dSODIxwoj9rnYNMCyBJq0pTGaON3OUX
22YRKOqAhWL7+t+ZYpAE0RxHPA5Nw69wgI3/IBCmyYVWlUTtASLlSHDIXQ15hcpcAW/kMMAUVt/r
IUCXjl+jesGEQz3Lt1Z4nPQ/XClHSGAtI3OQiHYlisq4ki+oBpGeJhqEBPl6os6KybPtbBDpYerr
jSyyZe7VO7jG6Dm39b8zPEYXNBDA3VXnUEOpftL84675+B23XNYwU3CRiwar6KBje3QijVwtNAii
eKhdXwXCPUBZDTjvGnNHeM3pQjmFqcebkhvqGCdIYCSI+bscxdBhP3lnqv74NvlFbqJ6x0afrevE
s2XTp13sA3RNT5zdGST0g4QIC4jlFgAyV4JVwjAZ/8IzVkKLZVVoPkmea9BPJp61ryy5+YIvwlpe
YtwTW4q0Z+8JTWAUEF9e4kl9eWrU6PFtfa4qQgx84510tyd9BwxsV0cnGvnB+PHkod2i8d+12SHU
Z19SMZMZN9m12g7TJ/GGys/Dp2f3Cea7qh8ZJHEyptiSsbG78IPTX5BXHScIvpAwRqkQViE3R1pO
WCRJR8+iAWK0er4iKQPjMkKPqVgxT2Gt1d7DzumBMnM209VY29t5HiLpkpafsNBQRqZJZwtcPApq
OApabi6twOJlVeeNILfmBP/+i8rr8B15dzPt9MUqMJ3IqZaefF378UQZ2ktQUNOYf8z1pJvZgeih
lGcuj9xGU009Gc8BsPoxqB5y/L71d91nzkT7DkErQNMbda5B2D/o6JvDt1quPYqEVrLnk6fsm+ke
vqpJg4KEesKf+SjZ+0KyXJI+Wxmx8cE12blajbZZLzjQ+hOIeT5yst5m1eRcrIwWtka0xyM3CAG9
Rwfk8b16sGbo1118B0zl62sMlcmWGQwW0FyPPr9wqkgvTLJRUxD6WpkE1yziDGd+fT+Xa22d7uFR
PZJd3hNjYl1dt0fg1zgxscPIz9iFs0r6juaa9Fr9HtI06cZV3xzt2G1LSRM2BHg4DY8raWDdA3TK
pIOhmcHh4Vh2xHuR0teJ511XY34GGSkPVMyZcjXCkyC1vT3JAmHuJ0d/six9IK/L1vN9AL0qTr0t
bxX9qNROVIh1ppZiOP+6qqTSQ92j3JdJh1HPhnUIXKrPUmuvjsULtxN6POsfzdiUiTlfBtQk5NPJ
Id/p5JJ6VSoqxUJX1pDeuF0BCF6CLjY8HGh6T1ZT6HA0ZtQAKmfMIbGN65ukIQ3tUulNOE47D9r9
kjA8o50dG8PhIC3xO4Qjpm/vVS935KAC/kB0h8Y6pjww7I2T42Ypz8I2XdxlpSi/DieSbcigivyX
OntJ9vidY37eqBiOlX/Gf2iB3Cvij2M2YUr8Sw98ui6gdYEoYfEDi+QUb+q2dMJwKEJpZ9ZPldcJ
PBo9wH98ip5wYjSlvj/wh53ySrin5Ej+83N3X2Ii1hmK4ZtZatZ6fbV3nOZecZ6+Om7LP6cuAKBh
Kn9fS3vqiou/b0gNMNqZ5EHxHI01aVB9x+/Lgf2kvtgwUV1mIF5v092f3fLTodbeZha92JO1HH9N
4gQ81c+T6FGuicZiJwDLe8EMnYOcUPMKF/yXX28hYIh4IO0OjDDKSViBb9o1c2PjTO+/ck4ozXTW
g+psbmduXuSeDzz1cDDeKHRLAC6R/x89sRhkQPxVoTjF+qhXC/bhjeAzIxc41rCf/Ezo+jqVvWy2
pXQOhakk2neN7pouOzCsPEVrVDSioeC7nfjMkzh+xhrvBeZxGuNS0d4PBR0g0F3vc4MH+5kvUoZv
rLO4ABzp5HbLOjtHKoSKvtFBDcAjOblXnIR9pr1NxWh7o+i6OsRQPguK1c/gh7Kj00//XnXV4Q9j
3BXGdHarQMhXATSYTrSWCyY7NsUGxcP5zQ3S/wPywv5me+O/fo3hQoAx3Pql5g9GTgdy4bA4HCKe
lbG1259nU6lju8RtpUncYLX+jpIposCJek5x6P9XhpQLKO21HdtPy5cvWbHRHoU6A8PXhZS1Sego
5ghHlqMd51NmTD5g+tnKZlkcC2sMJjJWPA0RJnLMqERNWmc3pWGIzTLF5pD1INl+UNaAnhOCI+Np
Irb3ma1tQ6Ci7vvpwLIEyXGrNMFobyaW/yHJzdGezoySbub6adPml2rHS0ub6QYU96LOF6P5B105
QqWFwzvxEjnA4JL7tWYvvc/Ok6M6zCys9JqOPnkMMsb4UDY/+J7pgO1Hmyy4SI3eEJqOMMWXoElK
5smTw/SGEQjLtM+xdQlBfTFuzhqOQiyYG4SznHHFpLisF6FpCKPMLhS/FCXEeWUpuFH5XwbBaW5a
hocvq0dWhQFZFDEZwcbzkhjLodI7XLY/DAeX25XD6yHoywY80xHTtXDIlsZKMqVzTFbOyeV6v4pM
8l+nvbvDyIbuqniunslTrBo1zmkpDpUL5qSsrnQDbCrlVkkTbXurt9r8nHZCUKDXz/m83YP40xTt
NqbIQlan3u63xvqBS+yX1PPeuG1RB5AlrbYYmud/tXlsVdW85KHfDPzTtOXY/jmTVT5DaFK3mve4
PEXpr39TwRPslngwD91McQdtgTLE26RTVpAr6DAMPciyClZTGgp6HCkvubqca/OhmytO5y3JglfY
EdTigb63409kIOdustNLW2R2tbpVvAkfekRGfz83n/mWUXtLoyvvEL2GuGH3QcafW9n99kFe4J1Y
bupVK9wCs+KRa66kgI/y41FJyZLd9cojt6A9Y6L9OmczzcXgCTC5oY0yxK8luH2OwUmFp9JiOdg1
OAzgAH9tX6wpKcSY1SW13CGzvsryV2vBLW8oZ59TT1CxiSgs11X5PzL+alhw2RWCRBnHcn1o0Ltm
9NbIVayO6E9JBdvZtjfsss+DOBuzGCODztwomPDCfCBGZzbCXBaw2vObnEYOr0RCbCa5LT2NiPyA
JC+x7LmdwhH+JHcCZksZng+S0HdScDVxMjiI4dJLdOzks8ngiy4bSAjPivfzu8u1RhIOkMf9jb8d
GSz86jQ4FSaVq/PzFVdejkl9Y2xWlE5WY3eH/aDfS5IPtq0GCyoRaFi1gHgPkdZ0/6VMA0WlPvcw
BhR7ejQCRGyuMfaVAVgBkNz7Z4kLt1Km++iyyy2C7B3tsiUtFrtqSPutFGMsTeFRvBvQEhRRnhBm
HBl9CyCsbQIuK4w/JUB3FvPCNvYlts1t8IPUiTE33u4GRfHhphuzeP+THprZiJOuYbgszhrVB+U2
WIdMwOy8Mpqt7e43qEeNk/BLDyj55GdMzI6y9+NTinuB0HkIxXlb74fedp/I8gFNlkTvSDBRq0w0
gEgQH9EHSmjy1atEp/allNlVydDVjlb19MKttSKw9q3N2yqD3yryo7WrrrlqQaEFAxYGoskYtb9d
cqx3ycLujYvQJPgNt+9FxZSf26JmW4gte52rjxEppJub/+DkFJpuWbbJ6MqI/SfGGQM5QMHbsvfk
WBbyeas3SZRxz2wXcE7UjabqXxomovJF/cLbktHJ5f5sX09br3Od37MW45GVReMQsCo/5q4s/o1v
XzP1AXk/LZCDa0QX2k+VBm8qADZtT61E888Es6E5QVBQPIOmGnPaLysSDNu8IEYiUZIIEFf8jLLz
jxQku6H8U8Ed5tKSf7gk4YJmtGxBNUDPQGv/MRXgZWEO69f9O9I/vxns26fcUrekwpqfNUAKVKo6
Yo8175417jB0UQ26wNsfWxsU/rVIKFYK4X4aGPaoqq2gUxK7N7VKCSiewgJO9JTzx17YeAdbCChH
RiD046sdqFZbGHyFkxZZt2CUOfTyRp0lZDWJiTCtUyUU68WH0rnpKNYky4yPWblc0A9cui/bJpPh
KnpU/c0yf/4QxVbXkwfIB5SOrUwvRQWwofBWrVQaEmgkc4LiUNm73rzubbseG33Sp/LaU4Wr77ug
xcarP5porBMiP0L1rPbgMs2bA0iKp29Jb3RMCfeIIEwoNpcfxXPflNJBlS0c8EmxCqJ1gC3XJR1+
ql+H7MdKKrwTyNRMn48oZTtCJNDDtBOtg6aEhNYE+dJAEupcttNxfncbNEH7qY+4gU5Q9fy7gHtT
oEPeQJbviyKJ3l3DJdBnPDJuTb5pJbKWpk1WeSNRzFincDZCRpmZAcIem5YreyfAChYUjlpg4vQf
tUESpAJknKSHOhhQsA7h7m9cifqWPgGumK+1YS1hswZlO9ZIa/sAP9AqrF/nehwWh6yb7boCzoMg
/bJ8c2lVmx6LmHhSbwwcmnX+wmYggTO7KUPEIfeq+TYPaF74lNdh0Ag6WBxCY72I+Woml7xVJLB8
yAYBBrJ6n5Jq6UPV9SV2av/ywSLgZQfnUnQOHKT5LCSfotOQxvefPwTMGzwWDIqQ/HClUhIvUWuk
1m0LF3pPW0pSPnuIq+zdS2xwurPaza0PtZgxubQbBYmqZpD6L4M0iyEM5lmYl/QyuM8ODOyyBm7s
92WnBiOHRluaFfiGEmnArk585Wso7zrx6IuL51PdhVu3yxiY3fNFJnZaxEtG8vYSuPV8JALvbMlJ
Gqo3/EIg8yofLDMJbigfjQcCm3vY+4Wv7HXbScZnafdD3Duvg1fyyL/m5/vAZ2ejv64N+XUUkcqI
Fhr0MbodPp0ejsrw0DHc6FPDnEoR35Bfb+UAV2k1XjfBMLcHPD0KSfOmnr6pHUBMhiGtjYgVFQpK
Gqwd6GVeJIRSqlsZ29Ku57VooAhpmeNEIeFDNvnwUfMgSqqTjkgsN9bi+ExKy4CZR2FEu3EwF9YP
6kxB3Inbk5aUSCH1Pgk4F4gspQEh2sWRgNtUuFQ1pltG78Q47mpDvRm6nkhN0jdoLRPOkDsxwO78
d1iG94K21JI5EqrwcoMIBwq7GFUUthCvu/o9I5H5aFogrDTMgiKRvhD+Bxx9XVZihkRs7jdzBRM/
+MpBXtCxLcdLlYFeSgfu/SZzNFD0pTLMXsa8J0C0i78yvy7M/+MYvqMchZD+Fttqbot0YgjL+vta
6G/drPEg3JfVkol71Z6fyKB6FaHQiLiEaL8eYGicGBMHIWgZTfowh5KVLy+Yg5HF1aD8I1Mw4AoS
J1MAxuCAkrF9GNwNGO4Eg7Zd5DDQgKgu2F7F5BsOyMmXiOCx7Eme2y/MCqErN0itcaupcwyZqH+g
L2Zj9t1s8VOFtY+nbcFLg1OPYkTzqcMGGoAqVYk1mbuKdQEstQ1t1yfnCsFptUyk/88mj5kPjvOn
kC5KWGeEI7jU2hgYQrUU93ypbPdPYYc8rY2Syy8IRgtBDidB5OkXb4TulNg1KUvdvVM8DJXu5Nva
siJPCPdmahbECuojrZ+tzlJUzm45AKzThCcPgWr1YB+NzHcEeFznw+opS1W/FtvjWpwdaB5W88q3
j4Yb7nnW/cFDqoBL2TvbA2o2DMXBZy010/rORWLRbzY0UN2iEp30T7CM63i0OKqyswLw0OstLHw/
laGGb5733MTS9emQP183Y80yEDR4VRn6PKrbaeNIfCxSezb6CXTBEDNPTlG5Nd9e8NCTJQkSOKln
Ul8w2sz5/iAPdn3xVTljPNvd+ExqtF57XYtUnW2JTTh58FkNv86DM+k2LFql0qb+zsT4D1m388/n
1kqRONU0dfxFnLoCZzgHxl/zYJiPYQFeDVaouY0RKaW1N22mqaiTjsa1aouMCWU3sQpoEVPNl9xG
WiD6UTw7/pY37zUOxb8lEPn0zNS/KdVQduXNt7T+uTmgZlhA3PyIQXDCcOb4O5+q/UI3lOj5m9oO
wUEmQxqOh+QuT2u5g/ARjoZv8+q+IUUCYr5/3cI/v/E/0M3GKKR3ZqvcTUL+hp3xvrTWzn6AaHtw
UnAgfzZ/c5IKtyYPaRlUaoVALLkZSIIBGZ/Xi3WiWl7lJTUfAQyhi6qf3UV0KQAkOc8zZYaKnobQ
ymLGScwZgo4pd3ZG1/FzSKax2YEPwjwriILT42Jls0zLd/xKl4uI3TBNESJo7EkgilPncExe+Z1O
ZxjGypkwhMozoKW41uoB6Ag38Gi+OsXRNNA1mAkjXLgtdagA6RZKH56sqM5azYhDM+bdc3lwPrlB
fN+kRwWKUaWE+xC+9C5Zw9CqvN0PsZutxfMVbPDenAai9ToiRAlsXfIQ5rIwyqRa5I3HfBSOelUk
1To17QTDk3YQMHbL2CziyY9tSbbnJwjjsXGCal58jqRd+G/ZqQDfg6i11xJ+4fyjiEcX+tOjcU+h
FF+hLZAo/NZbSICq8NK+kEjTNsG9lqV6Pb23Ou0X+/isV7qgxgZ5Sydk3797BtAamrZEIj/hjcZj
MnEJYSYOSHK1Zl6ICLaCyoR5OvgG8MXVZmanD918tS+dVytk/Cnjy7a81aXfUZanYYF6XOS8reEA
BLFpWvN0yP9zlmtIChu/94Zkp7dZUnoN+SNBm8sU91wQn8Ua7WqRnMf2yhLyofABUv1nObPD2J7I
a3bOpSLjjmYtffKsqZvQQhxfjqA+pDHiqxdASFbK6oRysCe3dAKAKMZMN9GMap2Yat+yItJahgT3
VlHPWGF5KIHoZlspNReS+J268bwW+xL5l9hUS3LN0dNtFzm6C6t8sgCrl7oxBjSc7mZeX5bbwrmr
kcX3iTOOcj3mst8dqqP/kEDXsIPOBrUR4s8ulyuzOn1CTUp1L3H3H3hj+juJ23SwQdEdZYE75V0c
MYXayF4bc+ydJQAUmPT/JHQ48jrm90n4DpdG4NWx2i+GrLkm2/3mZsFToOzTptonVAeOxKr2r5gJ
bWZg7rvJSyynq6MyrPPDClTsAMr8JflQm0z1l8ZL80cHPcY9AMH7QUQQaNMNCPaLuOR8C1jOJdvm
+Gd5Huldoa/d2CJ51KRwvDpUZ0wFKNq2EaXC3qn1hxuqaR/nukovkqXExKMZ8T2chi2vD8uSO8xl
I+rOK/rnNStVgswIweFKa54Z5CxURVdEvABT7PGxtHAtx6iTHAZL/+0M4U4PKYtoJSpohrqFf8D6
WM8k4e53EloRb0jVQaWg3mle/ufayZIXlC9e0ZKLY02QFp0aSWMLgzwKr+epfeRYjEV5+DYjI5gp
QtVpA0NR51sadDegpvwMELh1qKm63Dph5+qEcYVUsxK8rVsiRj4XCRDXj84ecIoCywVZHlb+y8GW
Pv/RX77ZKMUOde59tkbAs0F9XogTRjTKcnIauLswxf8Lf2D6dIjDCOgraKDg1kxUAhQojr4OF1pd
hvEAJQU3LXhmPuRhxWhIQPFtWshxJYm9sBq8/xcvScv9ZoK4azNGOfGGQQLNjckk32fYqkp/gFxW
e40gGwJ+gXggcdgwgB81qB7HRnNpiA7K9+SOAgvwlypvO0d9BseYHuLiNeoyds78D+Ws4AgUV8fl
FJSPP65VD1jMyRm70x87l/L40oA0Jp2LPU+MFdll0do9wy6NEiKRwbTMzVQF/V1dlHDKON3LQrI6
BYsxzzIYUqX1McjB/AXpWO/Kcam1P4r5+Qq2Ba+cmcRhLTj8I32lLiAfO9fgNeOI3WswN1BPsvSY
XNoAtI92eZLDPOTf/Dat3X2x0OR65ZRlbOQzAY6cgL/7gr5f29OxkhHJGEW2h7mM8VyI5kLY18B/
pDAPhOBZGuEeAQXQxEEj5l8Nd7ow5I7d99b20HkYUYL5jDw6ihNKvUEHzTreS0FxnI63q6c0QVtW
QJJSXj8S7Fp7Zr9khbiAL4P7X5up4V8QXfVYVTAE8q1vz/S9KUH2dnoDymhyrsMxIcFVj/AIgtdl
PjgFC35neOeGccpwMmAiU5Ule4NIH6rqiRvqXyw+6F770IK93+fZYg4a8rdgZIaFbWSDvZqn1C8R
rYrY2IY5jlpeQdTjiI5kl6FVnaLpmL9OjXGMpEq8qsw6eC4ysip6foyQH9vS5n78ri39BOh7PKXS
nUoOXT1nnJvVsAPo+zX+fXgay9vsmWsSI4PYCdAYoPwEKvBJK2ZoN4GMlC77g4S5OlAZBMZu5x6v
C2AeU00j1qqdBVl+lV7TK+TDR5lWOcYSnnFNrIEfDPAIT9RpEEI+BvvY83VObaMR22V1ZFGezhQO
dUwjf3ShBDZt/EzN8VabNj29LXRj8wDZaF9XnmXU/In/GndVDdTBoFnT2JHGsyoVYgcCHAO8NBzn
Xm+UGqXD05EhhXoVAuVXiq14WZ5QHWBZgScmEzRZqYNHSTSfQXJioqV+DbTpVSceTsqoGR9q4esW
Z8gGKzvlICFmoogYk8zqXAF3+GI5XS9BgW/s8NwnKQSrFzVttkOnZT9fbVAd28LzIwB5PTYZjsEz
KwWGbJ2dTxKO/5BPOIqrxV1bW9QUEIG36tkXMSwH9SB7o+4qoNyi5XalIXNR8tOGL8phG67bFX49
c5gO3Gzn+8reLsdKsLAWbPoBwCpvJuStYI3ju4Nfj1/SCT7D+Hhgr5lt4F4IIAu/QQwDgiB9GJRj
BgYqLv6gTj5YXQzttbpkW0Br+hzmk0b5r2jmXHRO+SFfk7+lb7kLBnkd0jlz8oMNIYc68j1TPoBp
nQAgBmzIhUPBBHGx9kBSUm33lMMZa9RLsTGN1NpNIt1QaEbkv1iOUV/OfDbI5MCZqCopOyUjgmt2
hsHLKbby+aiVXGXfsoJhQTsYZuyCpUG1pIp27dAL1kXLyUsbv0xYRGKkYNRh0THt5MPpKYmPUpmf
1jyUWWQbU+Efd7MMDbJllLoFSG8uFwH9L8IMSPw88ZwvhQH7OFTCXxLvLcswUhjmpNufOjxQT8Ny
cOHTI3gN6T/nxCYC+WHyFRAWswbrDs3WtrvIOrf0B8bjm4va2xuB3MZKgm2lH1X7G+RTVcIVo8QS
gYH4CuXkazWbWsKHv3UgSdoUGxQoVV89k+lUHIwIF5dN6AKqWKhZuZRvgc0YqhGRwExTliMfJNmz
GIuTMHRpvIYGIZLK92t2IjE661VjPQc/osntVBAiQPUfGtnSkUinOxORb1HhCSg9m0Dabi0NDi3h
X3LKRmc0/euZPb55DZDAPOE7ZQbjOpg7LPD9NrF5UAc4JoNt7sCyp/NmqTOAb7zIfZtcHXDO2KmF
SN0Zl35P/ILrU7z8VRRt4X1keT5WLOxD94YCBw9gg/1KsU1LI6J3fwKa8iGHRqgTVmcsMMvtPh5J
EVUR0VtZz7rN9gLJneuY9oLPo1UpY9kp1ua5cLxSaXlZNIw27j+75YoacUl2NqAmlW/1JdqgE/JX
D8vfdi4F0DqcqxQCZPO6TN14bRVSMxzFtI/4GqH6lv2Z/RVwGdpUMLN0ZbaAGHHPwbFPGOhkNTEa
enlsYX+O1VnyrR3bQoUo1vLQaxne8JDqqVRXb5pwHX15sG6sw7ma+4JCQzFXBiLFxU8KsQLDbqwZ
ItYEJoPGYQPs7wXfXYqsXqvfspJ2RhR+woT9tXaw2x3D6yyU8N8w4Y3NUSUvcDpZ3F0EyilLfb2s
FHKfujhNfJsEyVufur/2FRX7EVBVAKaBML39iSCMqrMv5Djxy4xN1JBoXtlP6qO+HscpJ3UDGjbJ
Ze/dymbOrK5Md4ucbt+R08FiT4T51cNoWL5U9LCz54Lm6TXvVgZNLacL8BA+OZ8fvUHxZ+iXqUIR
M0qzrM4dsK1TaIoCRBXgVeaOMQUFEkT/y94GS9ff85KcqW8mx4C7hZCFEes0iMuDPCjSbdklbJBg
ytIgiwsa3Y8hiopyZfofQn/JgBwY0YADnHiQGciv7RBEuJMT2KhT0V+Hyxp5PzVe+BXH2NUB4r87
drIntESMy6ZI/zaPYu8QXwrIFHxafiWEN9nZH4BzymC15R4hQOy1/tBnGPf4hng25AExpbsHX5tb
OaTptyZi0dcrMkb1DLSwR9RydqbxPZSPLUH3gLEsv81Xnv7J3tXIwtOV6Hd/H89DeNt8K0crsa5t
P32+uaB0ZOh7anN3HJ8KrDS5xF3Lq0UObrmuA72OTIHCp2qFJnVgDpxC+t44Jd2cXm/YvmRatQhq
9fg/Ykik3sQf6WqyRSOTs4+wrHLT/8rtm/ymq4AKnvLFYt4VE7szxnMityBf118QMM5e47LrspLD
iKKwXbiDBfQmx6JoYZUFag7wnUps9ouKkhmm0l86jm1sf5FctmsXvzYKlMMwxr5+8i8v/dxseMg8
f/W0tMskqwgyJF7P6M5Rl0eBQKAE/B6pBb7Fxqaqn8rprtVSsuLSq7+ENrHP2T1YJMlfm6v0aTwI
y1+Oa6QQv3zvqloD78yULGgPun9K53D7vJDiJUWrGYZS8zLF6DM4JzFuw+P201EH1D2jpwjGQQZ5
7hJvMRUTlfzzX95iDpL1yO9CfA8Xc2I4kc9g1vV796l4SNKONa+s3QusbApPfIBh0HCt/EGDrhU5
RojXOEmtVT+gEFtuBR+DbTbN8vQyTuklQN4p1XDXMB6fDEsy2hfEOshuLf109kopah13+ElDa0Tr
vOowUGaAS1BVCZVMuB075CMv7jurWmaIPA1dfUI1ieFpocIdmJSkQ0shZ1i+da3F23h886tDBk5a
xzC+AVSBUcP6RELVnmqVUffRBiV74SY0Tj8UKz2P5tLn5aS8KLEtxGs7JPmxHesD0jsSrMh0lw4z
8MT+IfA+8lTZyRzNVv9t1TEFEWvufh8n/EUthjxCZHEa3unmnYIO+GWUQzs2w23GoYsnQ0/lXms+
I4AvAtcemQ1cMHZy7O6zGN/zACvmDv/B8nFSy7fJJvdGUZdvtEePrPM6/EOEpIwSOxMNsKwUlkhH
LydTaCaifZgarvoJ71CyS7nraxz5u754vpMUrDBFJNVZ1bTxBRyH/f6Dc5rO1VpjYYluIjQfjK64
8neEGyQ1JbpVBFLdKzEuUNbBhtYEEWfwRtB04iDSbU5MyoGQP2gHGLBwMBWO6N1Pk2mId9wNbsHo
Zo0Ejqnl6XlDlDDRo4F4oa/N1i4ec/iBYNpm1QyjjgM9OjJgwr9gTLN2BALu+TAu0kFrWsFU7qE9
KFgiuVhI6eFH6ascSwmvo7Q1hslBMIIgz8EUCnc7YZnVvBNMphfUvBotsjDNvnpEC9+3I7wD0xcj
nltJk+7MRQ4DGNC+iEk90BcmHo9fJy9wjgNDHYOm7ysc4QUZ3vSRvvBnYa0syq9PwkSYQoKbDMXp
R1JwjpYVnxTR1pSVFqzgfbfyQ15mfkuXYT74m/Ut/jMeIL0F6TMFUs3CAqPh8Z9pqi5i1VrPZ8Hq
/b0w0alIH/SsRjh5R8l6rNYtz+GjEup5lfZWHFlVka+IumtUn51QnROFlVyJpg9VBxvA9OkBeRyc
S8L86pbr3ZrBM94C6rKemZAIZ8n/htbZBHZSJawREYIclcP4RcNjvVfuJHfgCNfT5E9rTLiOlqKv
/Gw9bS20s2uGzH6c08UlZ96e06zi+m2Kb1K1lcrO9F/ahocSrbnnksvsWXuTwd8gM8Pd0D2YbRPa
esJIBldyOqLOACngReKIjmmu0vsALCBzM7cJ2HvezLdgYO/asPVVT9OUchqdoE0FisBnv19fKFQ0
DUDqBpcn89mbFK2PFs7U+WIw1cdTUcpt+baEMI9cyr16glY2Sk5HsTqHr8xxeV/VdhMqNzqFqT1t
Iexby7ZIG3rYaGOhX65aqc5cdHyrzsVRYiOJShj14RpUFgCzcW7VjJ55zchcGv6aubDUWTHUic2Q
MhFZsjXCIb8Va80WD3kvHXLSB00R9GYU4b4DnWhslzjRaRZTyt9kQGiU/rJvS40W9txOSy5sl0yL
hs+W08kAnm8NeEBA0HXfWHyW2J/zXvVO5/Z8S1a2SrTBmLSW5MZySTgv2zyCLwUgTt7GIfL4vt4r
7sSB67rGs+kG4AKC/JyzMSoHMSDjGyVYSv81yJwlh9/9ECLIvXxkewC99vtRwpbiW6drAnr8fOzf
/4VVUKar5Yri+40fOEAmN1P1Ly1nXODkoekZNZfZibRTXZL8w1cedVsPS7xjWr7ZmPtzPYk7w5R8
DzIikpcrOVAQep2oTNXAgRJnCA5iZx8Lx6sVirPiUXXsTIjO0RD2yh3svT22GLOAKSTfU8iGcMOz
CerGqjZNXKpasJq1fl3ibai1szj0EuCTp3Zcgvfy8MGAGPONXbtbNcYk2FecMoPtDrVOqiv7aTal
10XFVnQeRjv7ikLbQQ7oXHY6h6Sb4LcK8wvUGA6DpmuzO2WcQvcObQDucTL52T5Yd7g2muDysG4Z
xZsyCRgZtCPmA0iaR5l8jlzdtSrAY1SCoelEx//pQGBLLGHXiONEhhPR0ZdMFS+Hp6CZTGj18iNS
G9lyQ7iJ6nYg24XchbnKUnvCQHK8Y5CP5euR035gq54c71Hx2GUKC5DbXGXdEBEfvUdvRmAPr7Gs
lxzu96BNy0OjVXI7W1FWSHB8ODYKt3SLR5LS1W7QjqhKEC7Oo4OdAtiU/wShM6KsSRZbwLlTW2PU
m4UBr/ZGMZ2EfRFp6XaM1XgQKel90TGPtxsW/Q44RRDcJV0t0uZU6nwPTKA8ocNBACPk7XxSSFRJ
oeU/J+/YygTrc/gGHRttjAwA6qOapxo6sQolO9R5pwxeNqc2l4ccXfy6QVwFYgIonEiXdwca9SDK
L6Z+VuPlAHZlkUQVIysnC9Trlr5N2lO5fQeiJK5vh6/FcN4egZXFqIY7InEVwp/4L+rE0AtcBv2+
49cOcW4OImaktXmAWnmf8aCF2VTLAjLZy/QKf8SsUStEeGyAmBQFdT5yFhwN7VF26Dk7R52DOnLc
2kbQLjXQOP2Xz36FAtkz4iY2BmZ1x3Z2exDTu7vmGjjSHKzWO3/nZSa7A99JgG4Oi0bdveik8fhr
3R23j+EccBWIKowI7yB2a4demD8n5uB5FlsU7Ikn++OZJCy8olEoFBM697rJI+mQogYAFiZcSBXr
h4a5PMsqt79kctR2jIAZDptVM8DgkfzzQXqrSq8Qp4wX/vg15Piq3PXT+ds7m0LjQcrWn1ywazbW
RGI+/FlASSAVLdw76Z3ifd37FUSTcTf5gzc07MzLGAkWhEBqs+T9yKbD2Mo0R2CYWzxl9K2KtNWG
u6QjWznhK7H42WZKTZpAFzr2UmnUatyUc+iozevAJTApNoxDlHgc0U60mbYMCvB8wvclZ0BFKRmL
IRfrvXQ9bxfC0xjPlj1OdxqIsIH2E8j2zT2kTpM+mfIFhOYTHqvGjn2+cIvUFo1xf55S5Dy8CXJ+
zKwNBP3x9x1G9lUDAMHINQ3NNBpYjPdjScPYsr10KWf1nV/DMnOHlY+hbeYsLlWlDOmw7Haw2W6r
TaiDcrPnt9taUy1J9z10YynMLYPizoH50LaYCA4T7nvhVZjcMoeLvXKjRwN6Fqqf0hASB+A+9ccC
OMrIWT73e5gyQ9bJOc1iW/Fd4+ya6tvmqZIEyeXVD1ZC+1CqiRorApLDkLmGkNjBpxMaE536nO5T
HPwO2hP9aMVjx+4i8nkskqSWtb3mPFT03/wmU75rRwLYwmMymrxSrQxc3jVESCv2ms+uZkYb9BwF
cnaikByIO+ODtI+UZuXwarM4zUmYqItRvHITBPUrWpf4uSs4ZghqNQWqYPE7ZP3dWkUjfZ1Y9tTQ
z38qSA565VK/sNlOK576Bl9cjqsp/kgi1Rv16PK0jBYO54dMS8qODHn7VzZ3o39aNBQlYDXB9wgh
Iu4OiyLwFnloxWEQ8rzhleoZkopoAvkPlhWoaItzbcdMW3R/FxCr9H2umbK49cXpoB1q7ftZSMx+
Xj7AH760ABvJI3KvN6Qckss/4tbHLsESLYutwkbfv/kTt2O6LL3xf8Wl8Z2e8v2VxFGSPWFnhchX
s9JUqjW1xvy3SFDDqn9sL6se2McVcgznUnPEpoLyyKa+/OBSgMt4m+FaxmaagjtsYW+FLJZRhXyn
ewP6jNf91aOtnDLd7lsDs0I6+Cjni9ldWbZH41rbu8GLQHmhflynY0OZILLQsB9zmJEvzQ3oDnSL
pQDJwlbaRSS8i+WIi1tA6vOPh1pulugGJW7Kz4NfF7Z7G3GfTSzwI2epT7WuWhIdBehL0XlIA7lu
gjp3X1L4yT1WDo+79IUY4dQ+d7C4cfQOyCiqGeeeio/0+8rMVEbo/G/ppUxaHOQ5pqEjGJdVaY8f
UgSPJLX1kEsvbIcVf2NOywnL5Yjbd28BGzet55bfQq7AyyciUYzXCncsA/j643pNoQuBaIGYzAfJ
+fM2MpUS4km2l60MAWE9Hf0bxIjP57Z5hcTIOvT9jLcDjeh0fT79cs3R2FPE5lGUHo4mhxDE/RpC
lxWzQQWjA1BPYCLmCYzoPxNj3pRzBNG1kSjb+XBFZrLTnZt2P/V/i9LxDJJzoaYIit57cQ5/Y8CM
+JM9/omvCGCH+Wki8TVlMgs/Kn8Oxh5M09B6eYFh5aOyv3dUagvTxAR2Rx7mwWqlqI5XIg3FxiZ6
LtH9YZYglOThEBLQoiTe1KSNviWjavskEZTdlIWXLj+jfnUMzQcc4jdm8q/bF6bcYZeUhN7q9v43
ARtiN4W7KA2YZC+kY37rhfEAGpMCjeNNH5TOMF+Zqe0+hgTI1hmVlUOcc0woQlg5FeRlGVLUC71o
G6or5Q/tt5tD97BOh36uOyVA8ZYjHxXwhREXIuP74AeuXC6+MxGT43le3hrltpwePC2m9ltjQ/93
JEjO8WpoK0ZAIyUV8o74joqFKV/8ws3T+k62QrfJvIuOCn8XJUcjh5ZUgdpeXxeIGfU+op5O+jeh
bZqCL+wF8ub9F5mnJQN3bRx6Yuwc8wKJWjZ8D9M2b1LnZUe9Cw7nMO846whUTS7BsvAuX5DNjBDk
64nE4fu+IZT4g5j1pnZdo7XLJ3vemnfdFKXWKLlNAgp0/pCvfxo/bo9hm6JCeJkbdAa6t21JzoRy
zUbQdSuHe1shK4Hmq2Ge2plAWmuRk5udfy5Q6i1SsA+NbN1GZq6puyIV1HUDPRi421Cr2PsN+nr+
oLlWuwCNxr5DJpJVkjo09yxfhfzNaDmrW5vU8NtAEnDdrRm1o56lFSiaAZ0kmgUU31sgCg7wVJaw
fcuEZryFWMsM9UAyNxF5uGH811V1zQxV2W4Yoqfpq9UIp65udHzCX/lVoU9HT6pqgd5ZU/fuhPOh
KPNHas8ZsejF5ywDCjZKskJckqJOnxz4JwcMdn4K3nDUbD8aM3uzw5ebwZ9QlDDbWfG/mqmWtHji
jSxlTWG73cqPmMvQZB6LeBatupucwLcd1n1QNz/cVfyiSJdnbM8SXYseDUVQ3tBeU4YFKjiUwkQU
OKpAOsn00KRANIkR0IsnEUW3Dd200cjU6C1Ir0NUxrk+W60DyeZFdW//FWMcsU2UbDTINCjeIfKn
yVUTjawNW2lsVxRAvDwA2IZEl3E8YslMyCXizpWoSOG3TdwMRN/KLLQhn59SCDvBSBqusqteuxY8
QsL14WTHa8g0SJvJCjjoQCL1PUbBumXVe+dv7ol3F69efw//JEVu+f/digIMJCFNmH/8qiF0Npoa
FFwRmww/gLmnWDiXWijGI2vAe/uOrnbkXO4LUOtXI0RfGRx/mm/7yhll6A4mFub/sRINbCb5E5Z2
bYasqxf8jPqMm6jmjmVyL/nIH9W1MSN3KiXj3RTerHNfH3/8tUVAdrD7TKyenBt9TVps2VnIbPhg
VZCNeYAdEm3Z4LLNHnvZ9qU3NMvo3KLv+CtsaB+k32PwYE7VZhJpMgtjGmI54W7jzlSoAPFHL4jU
77PzBI18YIwNzC9plB4SdjK/hldW/XAC3PDsqAFP6E25fVCzL1kRsxNWTtVc2GVKN1MUqmN5kCOf
mmEdTVkTvBbQNofiO574kDtoErvYWMU5vsvUh7HhdfKDWAyJPRlwoyiIrR3vWJR3zJfl+nQjvr4x
xEPbXgAC2vZDfbri9K14kqY1SVwMMaum7b0r3uBFYg86CnKEKkRwr7oFbe9oWxJLL4ELRYpCEpvl
vcmxrxo86gtRebHJ2oLo8TwinaYpD/iik4gcWBrVXPsr54H33d9AvCif2qRb2eEdGvkt+UyEOqvB
qovWAiOKqHyHn4JmNU2wpwYSPmj2Y7lj8SIjHM2uI2uJQTTWTu1lO8ezhoqXmsCOPV/YLpSCqzTi
I+e/r+b64txw8CYxd17z8xOAacq4W3nrDxiCuWeqKOMcpJ4GNpKEmNWGMHZPJEJqovixA5TPWmMi
VgpYeiWl0BVBugwgjloS33oj2c5kdGI8rzsQ8IKNPgxBCefc6Q5WG/UShpYlGRM3fWGShXYaDoHj
+QcH1Hn9ZiViC2TZplYgXTHsaGUECIco9+NgOVSBDn7aNw7a1LdmswzhIY+b9r2afx4aRdd7+mu7
P1K8OEHBaBKrtmvZzoPOOYFo0u8kusuQdmYO2NdBymI0yiVzQMhdufJqPwuzEbJxl2depH834Ohx
T4xHHc044wZeq2L8Si4zj/Ul1lLywusDzPKE176ePRznW6A70K/8fuyq6dRN+RFaxFnqnOISD+8l
MopMXQAD2N3qfs6kR3p3OHpbv3YHrEl5xihGc73+08Q+NFrahzXFgmb0UF4j8tFHGB55no8KF8ov
RRg68HjgoHaRz6igEDAKTQ/t/Kq1WaeNP1she7xzxkX1M/QNAL2gC+E7IM/M/Zx7R7RCQnPPwY0e
Ma/GnMGIcIbb/T4hAS59/fxd+k4r5eTYa1mTbU4KOZdgWRa+52W4/2uvKaW+4w8KhKTxC/zvbg9I
tbizUa9x5IeW1q2jHByKKhs2Yzc03Vu81uGuusA6Spwoy9uM7QioqIfyuZnJj1MA+Ktptn+JMqeX
j2SXKnebRFMek3oxpFbi+sQH2hQnIFcP/scJmK2gk2HG5kaXkxnVT17Q6cRmTwQ7LmJHE0baDn3V
nLj57C2st1O4VqIP5lJwwPYg+PSW2IzB4pt7UxkkKCIq4Tw7L5qd3OLB1gK+CmX2pBoMtLtAHNIZ
PfSlAZXmlbc10IbiSyT2SmYzRZ2/dM2PFd4/hHf9j2WhMa5F5uTm0pRfs7CBoGNJKERBnbQ0DnXr
a+DmV2pYxSPPrW/4qsDfEjuxEjzcc06x1GsCz5zeVrKlaKsoJ4MhnXtS2ND9Y3yV4hKLJfZ+03eF
g04OKUOQEekEJtUMqntEd/pOZ/mGuq1uLIozz45iiHM2Ue0JhhZ/7V/BkYEX1ocV6e7adG55CuIx
05BugPvEYNSpXxDOLNquDqakw+FnX4JXi7Aj8fZrgixppX/lIDiuQF9OCjEbo0l5r9M2NHpKzZFV
M/D211MuULOEp1Iwvwgja7rCQvsnNuYlsw24yUP13SNLMbwGpXotViUgex4E/uGEmGNSHNVPloPY
ur+zgmA8L+6scp85U1pT2EAWGFFCqri8G0cd4bI6AoTaLn2HSvNgRnHY46YBYVgG3cbIuE5puldS
dD77t7g0vCocoCXksQpn2MKyp6Q94+Ue6OB3hGUGI3SkQIVr7r69o0vvTith/QSz0YhHyZoiCBLe
JRVSQF2BheEC4Booj+NCKiRhHqcnO4fycmScDMvniPMJv9nhDUOP7fxqCZud3/tzsT3MeCJtMPBA
mzyhY7gaq3FEVmjGK2Yhrf5OXLJBz34x1mgMaOA0OxZYfVgJBUU/j+H0BLO8H4035srNDIhIThjg
87+9GUgo5jBCGn7RC6tRdWaTmPwDwYLCISYC6ZGJUi6H3j0UKBwXIoRlEIskWpwMcGgB16xkJOpr
9/9DYOKYf+GXZyqcSwXtiOqHVZhXu8dzTe1GDFa16gP0ySzQ+Xe8tDGr9RfBxN1XUvu18MAqZp+H
tlQqrK3r43fPiB0HyzodN6wcnbDDZlwoOI+lXZ2bLvTtm8fYvDy/8j171mDKyIQRSvmGWrlO6v9J
v5hKKVhMU+Bzw8BrcbCkIkEyTZiMmiX4z3tcmMePMcyPxeXKGo2tH7S4fb5o3HxB9K4MW4bO1zvC
YwIDKBhZopjhy37mg92UeLOZQ4x6Z1JfSGfJnoDvh/xFDsjjD85/h2jZsZ9ZQq8fZlxrdaZl7MZ2
wvh2ehQ88RY89E/lFoA1AEnTXB8lu5TW773B6PdwU7aNT6slXXSOZeWMb9hfH+mCaQCoU3yN/vCT
HUZ/IxBrZqQTxoR0lIr9sDW+xefPgbLo5eT0DnXVhiJigiTjtrYdhgVZNhHujwXH4A0XapQkButv
wACOJuxipLSrd78IZfVOy1+0GiLr6wkFvEltV/bB3e8YurKJrc+x+0MSa/nfuwr8eNwz3+rQMUVC
JOh0wHolzMmu9bzVGI0Dai1FA/Z7XTyAawax5MZFmj7oJs5Rau2VQ3QG0RPEuez2g+Aj0AbaqvGJ
QTIHYyBu2pFi8CB6DbXaj0Vo8GM1ZaWiLYSTncn4Bl3NBzQQB6OYOUpLaKRg7vP74f9IxxmzM1OI
3j1IrOnB+qN5aryHjSHnOjstEOPVdwWsRGKI60UDXrEBv/wEobFEd9sQnFStxijcSr/dAf1a8qoj
N4Uw1H1SkYkJNY1Pw8IV0mIu0i4htTYs9WMyIPZRK6LagC6nE32U6qVOTQtpAal6EuhtXU6tePTH
YrAj++0DjW5GIefJqtlRyQA7ylhWFFCw77d63NiMIqlgwd1Mw7HGWJMXIG2b00iuVn3DDpPttopg
qGrKtRGIYwVWu4WXlXF6Ypmjf+3mYSEtcrQiepPNLeX/m9KdWbqSqJ0eeT9md/zUhHo2Pu6s6UV5
qFjLznoNvidProspWdOQqB26OJdTvkfra3Eba57g5kvKASe1Gj41hM64cApLSVLVadD6BTlGSyMZ
7hkPyHo47KF15AA7jMPN62nr1G8KWQuQQxk9pIP2cNWgPMkylj9mOYBiRyx9SszdvLUs06ntxHna
GwHMSrODdz7dVOZQVOzRsBH+eFQ165/xvCUSdbf5SoO1e5UVVk07wRH0Sh0g9xVi2GQw8gXd5cT4
twAh678yqfU077D4dh1OAnO2Sn9JGc+mi5W9OTwFDNbbGPGk03oZKwwUBtDQlxry9qfQlThRhqV3
GJKqf4AQJkVF0yOMMtG1LiVlrO8vqA4sF2jMa41qJzjFDXTc+Ze9gSW2Jrjf8EuWP3aU2DBHjRnQ
0oSGUhlSQPtgT4HcHSuNY0TLHKxtLDIyqinkET8697nciRcnWAYuCLjFhJf+T1Ex936FXTbMj9l2
a8T8gYQqbxAfbVrrbLHPmRYN/y4gaK1ucirv4ek5VLFZaAY7zAw35Obpw9cZzIvrHXeHl8HPuLdN
60CYP8tEGqw2fdAQ7CWm8FFFL5PrQrLSekoms+t8KkdnQIynhqOQwBUssmN55Y05Via6QlH4i6GN
7/aydylYKCiN2CqV9QKXC1XEZ0MgjO03Z+9CVCUBXPHuMWP0dzDxb87CphsUOzHs+YeniNn6DwCm
mKrsmXLPYVcmvSI5f8/CfED1nBofBgxFTdLtincBoXhZijR6krM0EzAtXUrIfpej8YR9P8QwNbba
h2aR/hoEGkJmGmTFS60+tAnUkIvShCQhmyHFNA7y4wX7ljioV/BIzX6R9v9sgWjkS5o3scr7ssmI
ZjHD1OSpv6OSDD2+FqGibXt+Do28D9rcWaqnjziglmBnnYlWxz2O7KdyDRS2NvN14nnxeay3Nnt6
1EayrmjGjU7Qn1EMufDVcFl3+WZwr8zsgg3UYS83gMfJwSAPv9ckCnfbyfnpP6KHLiIFTFyssbiQ
emBWTHIPEtwowXMI3sId4ErArWUecklcKH9FtzkBGwKnclDXYmcK3oLSDeF9aU/EYpJacZlum+xB
IUb9o2ESk3Cog8iz8Wj7Spaws/fzVSakCza4HpI2mdg7dQVA9oZVXcCSFzY6NzwGQJzGJkSUF7+I
7GK5XyYC+osRtLAZGyrR/vmreggtXOQn+PwCv110HZwOYJYBeJbbnltGxgVRraONDtSt+GqWHJMP
GOlB1UmbyQUHcnagjJ5stiSoHVcHx+oTX7s7mOB2ugs+DTs+3h50AN9NLMSxOrNb3q7k57qXnWaf
IFAz9XIQjek7hbqL+cSwPHADrkxojaQWbkh7OnEe5T8Qdl02Uxm+2w9gjD0mZGHsb51AKiU92M5/
m/VqMGCbC5CM0/eFD1vhQ2LHjHX39IiPcwjKznWJPvBiV/E+fj7QpVX/NE3tVxI3nVvjslMriYHa
3dfazfOWMvnJG24kuMUPhdT3W3+NRRBp8eS5/CtAUSKkRBgK8oGPEZXRgc0BHhKqnKlRoS72Ki2z
HBWq7PVRxcPo3V2q7tjRFzWsAkbKeTr534ELH0WCFsLuZmMk4WCYSjzotWlkFvbT7OtAyKJQykL1
pWuqdz5q/5qwumK+MX+ub+IrKGsdn7BIkiGAyIPPSoYso+mn7MtHvUvVGt3ylXG0zEVM39UZoeDt
e8hMiMOyDwCZFFizcfMolB7Cl44SRoleHyWZsRadxAtRs+GBKePYJPhpm76HFTwHx5GAcJVEAf11
Dgs17rPq2xHRh31ybJZ0DD465kXGGKEXZojOzc/kH0YO1/o8hKEp5xqeCsNMkOOA86fbXs6KjNsm
+YRQjfXkSCPUviRmOZaU0g+yTO5tlyXPswqXY6ih8L9KHa3j2c2yPb0K9dPJK90voIwA296LX4v7
aTk5LNkmtY2224vZV04s3mpFgT4p3e+iOx2x0G0CdB2RN+tjIM8EmU7xb4k6ZfqTTcnBM3xZi21e
R5+EAj4uP8PhVzpohjq4diKxS2H0pQ5E0GLc2CetSbLsPsn26BFH2CZ9jVsRnmvGnXAxTzqUEYZv
X/dZnXIBmfUnyLe1ss1Lw0kK30PUKgPsDoxy3QgrJZnelJJxj4ciCJHSFkhOdXXzT/4D+TE5kizO
iYqIXySZWyI/DtoMZLymjH6AdjpwWenYuAvXbjjOFYzOkCub/Z0kMexnDIQvNs4IBjpJvWektw3D
6/cYz3AnW67oNuKLHAA+M/UsO24fH4ey4x28iCfr/kd7wLJvR8fPc+Z8YUnOdKWcPBo5pEhQJ1yW
crCRg1cSHjlbulgpK/sXTr42aChQAC1NxRpMkVh13AZaVi8Td7j6ZxK98Ek8+13AHFuVVRKnckNs
jqwkiaeMgXs/eY5okZP1hm2VQwTa0SixXPRGql+MMUkCDc5555pcPL6/h6YFpMmMM/8KFt3zGImG
wnUqQYQUEv4zXpZOeO9hdMLHP5fXoBbvTjywwBTeGFWnE3XfnF8e9V+amtOy/OQKOnKZtcMnpYn7
vqz3k0tbH+M1Jrb+mq9hL3cIMiknqKk9IV2JYntFty4hyMcndGDXS1hUcyux3qfKAb77N2td1O2h
u8nLSIj10kZTRRvOLN8FMVVARmIQKvUDC+K/6Ll9bczH+k+4Rh8GVAy1lmrGHJB+kzHClS2u160Q
tO/ag4G+EmBHRhmcvf5haz0FpIjpnW/+M8OQrSfnicCEg2KyHVEeSucZwK1pb9qN1lj3cIVOLfyF
wSKaS69WIi+c3l4JcYxNWaWUypLngsAK655Su+j3uI53tcFoYViwKoER62qC2vBJhZrpwM+98iY3
0HT/HTnSmQo0yzFFv0kKOtIle0FbFeTPYdqO3uLK0sVBPmmjV36j9JHHdtcwuOnP8dtKyqH676FR
BsC42BAhPdqVjveuiKhLkwjmDj2fLOF//zlffcy5duB1yA9ijuL8xRI6eiIxREtZODtItIiLvwNL
cIVn3OLJ1F2SSF4vU4NAyGeks44AjIIKalyO4G2Nw1ZMiAzKZUN3Lx6+PwsH7mAbeSWsleyw4yXQ
pnNGWVBoNbHFROG3Xl8JmK9WN2Det9AHtX/Cj5clcNxhWrlfvwOKAIW6fvev7rfg19lvyHFwd6Hd
vgSNqswsqhp6nL5VAF9oX9d43BuEcK2kcOnM6DQ1XEcf8EEw5T6Bi8CwTbf1Nc+vWBcXC+nDGjML
Bg46wOJwtn7lhJjLBbA3R21iepkRWCHUNj4grCa7vJaOMh2Th6wzd/EvSIBgOw5DSABkAN7S1tS5
4Qkd47oWtmuuReNwRpNqvwF5Jew/1FB2BM6PZ/UgkeOibofOOq40jHKESwm9oCXbc4caBX2n8GTb
hoh1zOrYBbY2856JPQrwXbK/fk1/tloH4kMaAMA0WY/YbhmYV2IS31/cfveqH+acUG+nK5Vbj/t5
i2Nc0ESa36slh2vSitqdv5S8oaUotxsCc5P6mdOj1nRZeqtxJyHwRNkgg3X3ELQQFZz+rdqEJIyH
wWsHqS+ylzFiBpqyxatSseG/80I5qB1TNDpvERLHL27wtW3e+X7v3bHtdpFiDEeQHF7vX+gEQLnu
f2fsEilocCvZNUZppn1dTtTNPEvsBd6Y+XigYlPsKDkzUwBsWUjeVMTpUa2HbwUIxYzu/b1wO6tp
X0og4jF0FUApuvR+3G1UTfFQgyJ1l4wdDgAd69SMjANWY/1UDBzorpVUVLrY0sivBGD2cYa98PJk
Cz1BU3A1PYxnxIkvO7QmzxPwljnzAMNrUoiQ+ojdolyD5tsUYGovK9ppR5lztDg8eGzcux2nISHX
/zZHgxKQoW71FD4ZfZiYEukXHdQtmclO8T7TOavVi9jaVHw0akK9SjDTDG19qiGU5MyomsdCGr0R
xPiUadgknqPskifbmJhlIluAo9oMMtb6+dPIirMNk/VDidpAMD501pAly/skTw7TFgz1rqbY3T2j
UG+gWjBURJGwYKUJuUqk+mYnJym1JDF8L1gJ1CRPzRQ703cpYHuw562gV/weFkKQMk1Lqh48Y3OC
8imXpohwjcUdSEHIpSRBjPWBQ4f6f9ii06/HI16HFUbGS1EnLHgEtcflWRqZPZO7uRwnJ7b/Okjy
SdzJebTPyT4jA/iIhr+eq8RwcwDatILiAy9hKrtDca9U96G8VaZNOzou+T9WCvbCWglN6CFmiLwF
B5wcF1jOppps7bNJVX1UfJ1eLlEaLRZkwM2Ljo2v3YhXHmSB+HQ6qwEZgBoL96IBslsEAI1SjaTK
Dv9EgcBvxxe9bgLE/o9lZpgcePWICkmQxgUmBui+QkNRhIu/RHcn36jfBBHjSJTnqKxYtkaWfA4Q
i27WK8xt2tkqisCJ6SpveCo733pXWKyRReDLhD538Y27L8M3brB7d8nkqs6hIz28C5i0Pfs4qAhY
RHbCn/roJ5lNdiCFfh9omM3ur8SDNVBU4j+BmfqeAde+u2jtzgrwMRVM6boE0wf5a2J5AtnMzaTu
pRV3i0MMElnC7OmaQJPvgx3xTRt53nySRiEm5gbaUPePtCFXOSBIIjzUpkqYKUhyYi5riLOB6s0G
tvhWcf75/i5ILyj6wuUta8Cd4fKalONSQRZTL1Im6lgYqNVOXg9TOZd+ZONXciMd81SNXTq4uklh
rHLP/mlkQHsqFMh82RH6iTH+kFGp3JutOM9SR0lu7Dij7QDmivZ3AAsKxSZVy7J7ogo3FuejFGY/
jum+jG9vd7icZqeqM1Tp2dsPDgYONgB+T44dph58XSNlsoNwGGk48igA6oFuPgz8FBOe+WPrcnPH
VcEfBW1id0GoaiF1QDEH3Ha32yiKPhzG4GoJXgkrrCldErZf1ENv8GUQ7Cuw552UBjXrWqnlO478
BZ3HhV/9mULBPLhmLhz6VH1TOoQKI5WF1t9uAScRMa8uzkEke6KolxIBk6+ne2s7k3liwN/5PC44
HvT02+SV1UrdNr72i9vGX2mcF6GPsGtScNAt9uI1WrCZn7YnrBYI4eit9YWRHKbAbnz/w6B/fKCe
ovu9cHzDBhN+UL4FgTJLlCNUGowdqVdUXs6J5AMC69c3djSTSOL7+HXfptQgQtbRYS5NmbQZ/xqE
MuBIqkNrzZ0A6RXyQQZxZhA/Ux6tX7IymQ4MhGhVeQPoGv6K2IgPKvq+XWdmYAnHAbOcYzv9CEze
oG8GB7H4udYrLqxR6uH9qHoxx+oTqdpja9r/9DK0feIc0JzIZHw4oqj/1xpdtNwZ1YlgEZaK0XaV
gMMfsbzWbFgCreEfYmZAWgY7EmoLjZAsCCnbNkOkq3sYt3+4USCuXCnQNUiBxWbMliXVH84d1BTT
exN8PXRC5DQVZvNrAU77SFXAqjNGJMaKHBvmBfWPu25OgkESffC1Y71iR541m1dzXaAw6FAJcQ4U
7WM1KQJ7mppuFEtKY+J8yLwb588u3vuNBoc/Uidom9+4iTwU3PqYiAdVltrJTzc4gDQWBzRJ8Rm8
KolQFZHcQU5woLNG1zCkIlw3Psf6Sc0zmQ+5aPVqJLLphZpG+Zudwy0i+zY3FeRj/Gt8sxOrFKze
lSdsj02iMK35367idUvXUg8toOHkydCu8n+iibuu7g/m64aAD8zYTdq+BDk6jpmgvvqCh/ZY6Uzh
Pl6wWWzMA3aZJD9G+3pCHxUuYHD0awKmifkD7dLaG3w8UYsru/064Dgo13LPTBIi5HJj2SZgP+18
UpKrwIM5jY5pBxXvV1ZNszcGjrXy3a56OL0nxsfn7XqGSyfQAXrB8x2YAr1Cq+QfArpgdcW2OWU3
kXa2/8vLc9yVFEDAWHObI4ZpsaMYwRfXX+LomNWqtiTxcCTr0Grs9vJqYZFkV7MH/X9CCOJmrZ1g
SnVmbJ90VlM6aatUPIiKVwlk2usZw0FtwzCyeakIgp6Kju+giMR5oGiJcJl/a0SB7dA+/V2RzEKl
JilGIbSml9eXOOoZisVmm4DD7P7WOzB3aPRJcDR1y9s2tXR5YW2KqrIDS8EY1zgya9nHAt8iPYk3
Rdh5HVe+xXZ8LiyW58sFcn4Oc5YopoAKNiu5FQXBEXfdwgAgPqnuhq+83tnef2MVvRz0FrZVK+Xt
hhqalC9FPBmMLq1xiO3Z1hW6I1MjweNMaTZvQCA1xzSMXOmzrpl4/FKxQfa2l/rVbgkhEcCWv7Fv
jD1Px5JPEiNKbvJx9fPElBQUxUYM4XTjPiUHarznqLOBy5Ecr0n0q9iDRYHfofMohIbS+Au8ONqT
T8X1GOGQqsFet2LMrT3du19S0NE91iGPFTGewf6Iibw9SfshtMfAffOu+znwONySp3sRqZQX/alN
jGzWQ85dUkY8JnyI6PEl6Y/OOykY0gAxT13SCeYMBmfkVF77C1aAUj1l7vEVuzZFy3AAEQDELiXd
892njtRwcHKlacjS3bYVWraNRGP5MTbNn9Ug1eJP7Kl7cy4mS0HIoBhE+LBGxjxDL124ArTRALcx
Tvj4derOaPorbVbDgrSfwXGyPL44r3jPIHtFQmozc9uOwPpHSMSo4U7PYjEq2OAoDgh/lbWu14/E
441c9EB2Tg3/WcJ/jx1Cg1JjXaXC5sqJ3zWyvQyuSQr3YD16mHVWwJ2qamkTS0RFDvMKLxGiugOX
Z2oWuP7gtTaUSLhOwXGiAaJ6FA/9c1AjXbUEoPeTpjYk3sjDinIbIz+g2lqUoRkv6lNqyLYBnpuA
P9O9uLiSWWlnUNArxNlqkilc85Xmwe/FVqdo3w+ULyZdnFyucnu1BIoeGba1f5KrTOZmYzlJUlvy
c1agid1O8nG8Nmi9GudWfYor7kIbjg6y4qArADwyEE/6PWRzROiOvxM9khbuIkiFoo/qKoVn8kGo
EqpoUdeYrsLFc/uJXtQJwX1EwWfGB2zcMMzWafqwja7nvLQ3IpOVwa0jmF8oICPlJ2yBBLZpoyeN
IxZjhaD0p3mNV3FCk2JF++1L2hDMB7/uDPY5LfII1mu/i8rbKRmMnWaE8mH2d/r8O2jGTEMDU/5t
RgQvcFo1GIv/eLwhWo0vi0TJFgkWtK3nSDclgy6Q3C4ghU0FRpbYtEJLsN2QFgEOnADlFluvKwaD
63rrN1d9LQE0n5MLMPX/F4gU1bLrGwSNNpXuUW/IjUq2KHZZC5oo0kUjfLl+r0XQde+Sf1WpxPz6
7qxui11HTOY3tkS4U70H4Tp70KCiH+vIHyxelt5pdZcko4Pc8Vhg6RwVUjMPCuFOB1/PpkthFrMM
ISxipyupvJzC7X7Z/swITWmdiaWskPDc+8JPNOY/4DpSmikBX67SsENrMaYo5149lOD3J5Xgbljx
0IcRNShOFm0hZDA1rGGn/a9a4TDZrJFQWZq2JC5wwMRQb87KgL35oVwgWGNQlje7krJMccnQVilV
Owsom87riQHLuLfGAZVMaDrEoE3OHXiLrH6NuYohtLPyTi9Dg4SppzRBsyfijku2GDatg1NzsHIg
HQSXUNx1rqsPD8Ht2+h2+D/ulljmAwTNc0gR+4WMeyVylm1RbFCA5YSdg/L0FPaBKlgvsthCIz0C
g7zRokCVb1EapdNKlu0OshrnG89RRs+3Iqb42bLxFksIG3STo3qIkkT0JqfMAWjiGWR3ZHYfFCpS
ntFCamAV9foVqz+y5geCqOCUDDNoNtDGSAxhyYOQowZSVCDQgdPXbnODumiDa2ej5fryw1cGkBYQ
nC2W/cNPI9GTMTPzmovrjNzA1Auvv8DsfryGauduaiM9YZ2K1I8P6ESKn6HGqwTxgrfAy1lU7747
dSPtS2zF7t0j0tMx7Awy8J1Vn2hHDYVh1FfNmiq8LVeC51l75XE3YFRfr4g/VYnnRgz9hFWTLTlg
xhJYpS87mpIb/liHY2HpDcwT6WQgaLsye5ueh0GrKMF2yDLN1K/NkCZYDHDksoyQST8WD/8vQ4N4
TssnG3Mo+lOXVFzyVjWyLjG+ehtp7p31ycy/OV1lQXrV/m55vz/l5IMZmjXFMqRK2tPf1UqPSwS1
ccNeODLQcYJJXXB08uylk2MzUwUjsAzQRnnXO0G7vPmf9Y+dpaqw1uLAYjHBp88V9wjgJfmnThq2
Q6uwOk0k7dwp6KVtWwVuWgsFqeMMp3LpvPSEl6rb6lgOkiNv5SJzA1dclzuxHFdy9DSB4wBzNdHI
rpg4AViTPHlohz4uvKtp0H2tSZJpyv8VRCYklAdKjAKQ1AZt27GqJrmO4gZ9NIA84gdnYjLK2HjJ
S3Zv2cgZP8mfbLYlAOyXsN0RB4LGWYITN41YCPtj3kCkzqnuXr8gF43p2HuCGH7HbEa82b6NxWa0
9QpWroikKjd6SPGa2WAWY89PvHvFM+Y/tpIjX4lXtMjCg/iBcLPOx3AfAiJmgjNt8bbZQvCabDXc
58KyDUksgqFV8ezZ0Uqc0lpBc8SeBTppSiiQFIYVU+J8yKC5HENc/k67oFKEbRnh9iC132CpVnbK
X88EPrNomZerrTB9op7O5WqnHirlZKmU1pQ4G4K2V9SnQU6ZiUgfpUiCysytQrcWwhtGI06dreVX
hLuj5AfOFZ12AJ0hQOCLiLatG1/hilPuHrRHZbxCk8hJZZ2Nm/dNTBbWkGH0IeAc8Y2dE2YMiyN9
lvao3DQQjqBnv2axx0GWNUaJFnKUW8PfTWaFY9toTAFyAsJUt7NnGM91i/pyFehEImqInHVjO7Xl
y4ecHRJJDGY+nIYAHylxj/5sJA8floO6d4QQBTdD0LcPdUUKpmXS7SuHJkjWrGH3HlptBIChGZ4e
st0P2Ozy5R+nLJbDSgxjqsV152wlQjc/qiOR3gQy5h1LQgISrv+ze6UNFaYmriYAlG3O1Y2V24iZ
7OcelKJz2j4pKfKKF6LJVTwlFHFhDsvXc6ccLI7lvxllc3q7lPfuM5GfOG9GfBnbrPxAebNAdLVK
wE6A+E6O/7M9z+1WoiaQK6z5WASAZcOijhZApfDt7nuN28fBvmnifxhtTHhNtCBDZMIRPD/lfXPw
eQGqW2XIk4idRmonwp4752f+Fc2yGAJ1KrFAXOXstffMqs707mTZzDChXV/wAEojJnM2o+QcYqhn
u+u+GNgNz5je0pU/lULdLGe3/DqRPB6KHfaPb724onIMnWRfHXTsBn3jKQ0jsD72vwEf/oaKso+F
jD1MQfh1uRxAzxC/OVyc9ySJjrLb0c1ayLjcw1FkwHT+Eneenyib22im75C+ZFVj5FH2uL6OI3Tl
x9OjZ8nz2EDvBIqJobAKtbFmtzMif2NX539YdF4KMDLN/oP+dkqWGv8sc4Lz3A262LtkSxs+xAy9
vt/++2zObd2lUH9OXo/jkYqt3u75jmhESm6z3Ktmn9R8UtwU4GCzswcSjrMOCPDt0wkniRY7jOgJ
azcynfzOSIudHXttEsyXNMJIYHQUr1EzCsUirS66Xo5019Tn3FaomczunvMmix/IrUnO37PVKe8q
Ni6nPmv1xcan1P78DcNjRArJFp5A/b94JiYAlpM+20kIEv44QiLE02QI+THqp6G9YgllSpaKqTCQ
Da8BOCLo3ggCTrLt0h8Hlk8bcn62e8PxzthIK9cSUK0781IuTYqOcUBKNE5ntF3KexNvfBKd+bGa
wQmsQOV/wDjuEdtqEJF/yFzOulchuB8yzSObCPt/XV7itLtweHYULov4VNAxmTuCD2zygUc/yXOF
Bk/eVdsqaD+55drfSSiqHrzXluzhUw2cKum4+LkPA1sGliNuSrHtEkXwPAIziDRYq720dQP87Bu9
3KSxjapE6U8Bn16jroByj2EzFBlv++qPuvetsXfAZXKYc1EKt3h47BQ4nvLrRc00kElx5jMbQAg+
OuMJg+7TSKy4OWxcYT/a+pmkcd9kOPIdkyh/K2EldjDL1P27U2CNLAJzr++Q3+XZ2KHmidUH9E96
CNi6gBtwZoSK7JrLcrooD+pqfLegLoCU3RcBuNz0QeJVMWf+Y3v5iUgpK3kjcrfJwmE09IljUWc4
Koqz9mRmuOKBUoKPX8G/5XbYV3g2GKZWaifE8kzj2EvIR82lSliuTOIYFOHiS/CDz87gBslWTrIO
GERGJaVd7Vr2K57swDSo05Xtic6OpYkd8YEpN+2oMkcP7Fg2/ng/LC2XulOre1C8MnXCKEtquR38
h9D2IZAcXZiFAlbKnE14D4GEq4qIduYhXXaI1Yz6PRi46BYxft2+gJfI1aSZ4vlwRy8vWCwKHQRC
LX5U7bCDwZSR7nBNp47QbGLXMG1GeylSZHtQ6JUk9S5DlvvBOKYB6L2a7oPyvWX0cXWYibJfs0F2
am8fYc5ejttIh7mS0NtogfYj70VOzSDJ04olu8CSFIoKO7AS8kDEHyQwfMQLw7Fxq9bfLomHWpPd
xH6TXjosnqFmcrsJ8uDr7iV2Vd5zPy3W5N+VBSqTPliJxpRmuMLDit8FQFhs4S9+94ZJC6lINjWO
zJ0ObxM9qapBcyqsPaFTt0lGQfmbRasVjOjQYBlzcrTo9i0i7eAK/Vfk3Jslr+xbY1Z9kA7qOybf
5RMjHCeWFUdCpt3IJBe7qILFqTT3egrfOblUI8o6QyJWHFTJZkdHcYE0kxb7YjM/U63pGC1HsISx
M+2YlnKOByST2bhsOIRz6flREibLslfTgMdUD6P5isNpcPjumndzrhe/uFMB4vzn2v9Nnz7tTYoc
lvWehfLib/04RLxNUj1Xbl3ONRenfhaqIZHVFRqiQmm6VZXRtirnpp1suPttxsl27H0md1gAVdwq
M8jNntswYbY9OLrFZxjxOQb/MLusLBIF+DVuPuHd9dAKRJGThD7Ujl57l/90hY2y6HVAo4lqLBFd
5krXtqCjBK6t35BPHculF8K1AYcAlcz2TaOh0afYubO5/m+UMZi56IiCt06jth9Y6Ni0aaThHZa4
zkPOmmzHFKolqISuxP50mr8NJ1POCdj2cudKPRVCWXjC9SFSfgrTL3XrKlG3zP6KfDI42D60rCqM
OznGtaDDv0Jv6cLgAJcxc5nc7TC6YTpBrePkTE5cejn4R6a+tQ1PBe7fmmLxgxouMlBF/nxlS7jU
OhXWdGHu7diPxHWxDJ8pOAaqLls6yRfNTracBuTJCCBuPPSSYgP+hR9LjZ5HbQ7U6LWij7xlxsRX
ewMvE5uFIk8/pmVR4OHTw5wa+ShExjDykmOPdiNjSzekUk09+Wnv8J6lwDUSaWkEIOdtCJhPwoTN
h9P/vo6pYAY9Cmm7OWSeR9viue/jE1ey67E648uo5MxqaF+SuIXhvDfZuCZEg//Rm3/bgeCx+mLU
KS53hv5+iTbDtRlznijKBSsSehQ8uifoqe0aZki2foCMJbSxHYVDWb7VHcKQB49rnWYbixnCQ5nu
MpNMF94KBoXOY0+6D8beB8/yKRHYa/7fZ+o4Mmq2x/Pj9lHUsZomxrRycR5Ccuul5k5Az502ES4o
IgzZNQxe6VY+YULi2WwYSzvb91TrUrfPyuisgIpFCinSygFtfxw4EF3MhSUKcQ5bORopomqYdEra
/Aabura/Tv9YNx//VJrk9+pVdPj4gOdsfzkmRRLBFswgoNPkNnVSvzGZoHNGVI+kAa0l6ae3oWBQ
HpGcdmkoEww9tOUvpQECTfi7N1h2rSdtp5UkS/5bS36suFAlCZPbE+Nei7W5A42dui7KhL4Zk9yq
DLhnhzr3AxgYcEtgCFvAceMvyG+BttzeV08OneGMl8dRtmX9kk2NbrO5D0IPLgzqxxENFWJlJ6KW
sB3FCoH53Vb3HhKA3dykPpwXRciGrLnCMGLMBxT8hpCNcx6/7drCOC9eXIg9EKkTgS/26i0GnOTV
VYGRxXU7TyihUQXE8aSKWNI2xFukDeWNrT/nqQOSLrP4sSRX3haDPeUm8DfNtl446L9zaVv5WldB
rHb89A2OoErY14+aMc7ve+EZdbIDOIud60rGy+o0WGVv4nGd3s++q1B9+Ko9Yh98F5EUoLoOoSyq
0hHIZ42fMABrJ5dgdOJKjYAKHR+uHJawQkoT9suxh1Bq0Syqz9mUKIbp9PpmI17G9FJJwdmYxAIO
TolZshIEsS8l/pzeLuZnRb9PVl3xB6ISJF2+mKC/zsuuKgMb3G9+M8bn+LlZ1rbe7iYipCaYmx2u
CgLFvefHdOg2Ys49jEX/6E8ohmB6oV5vdy3tC8OQHvmTlxQNmCncg/kCJ9klXkdSUbzPY2hs1J/S
EsZ5rPSb5paE8GYfVByekAR4ib7yDCOZOiF/UoCbZgwhIKa17oDrnq3+h0sK7M0pqdmfIBtplctn
c0un6m4fJsSGT6sAKOHgEMYBWb3GrWN4L+gwlWkaLWAs/t1x/KxBRlZVyjEG27ZKQ7xMgpMrjwMl
7yGRa+ziBCEFPXF0e4fyGmU8n10XzzQwYoAMidJoeksWUaHiqLrk7KGeUsWTj26VWL8bFxyyH1EW
mJmnL0qTHwxcXZwWuoS7ukZw6qvdJa4qPCtNxUJk9RhcKxwJNqvaHAZnm+1+93iTDueS0IzivLl6
q8WAGkPNKARepI4Tc0bVgudEv3nskf9MBemS8rPhTObepcEo1mIbGPIQMh8MXoEvBhVeKg387r+9
rwXJT9RtACI9xtzG2P8GQrXttrLTeEM52Vq8rglEmBPdf7z8Jx3xACp2aN2HIzb8I3v3ilEoHFaK
Je0c+8pI6b+yzc+FfmFAKB6RFPlwAH3L3UHKjYBSTx1yEtMZ/je9IF8aisT/SZ5U700QNL3Ck5II
YmQ1idiZERF340qujYmmlyxoa3/xMDJyPvoc5nJjIK4C5jDM5y5fZTP208/FxMfFFhl6teUR0nMy
KgLSQ6JPzod55FA9lu8RbHTnuFuQ6+CaelBLS7Bz++9/8IOcA9GAHQ1jxFur6XnbS6ruJeSIY7eX
62YtoTY4qtTuj2jiP8BWfQiA+PL339LYyFN9/oJSp+zG683xqIyvdRtY0+qyJj1enfESVq3J8Kp9
yLZzlDwSuUNWKEN0HlqOff2EImihKhx/wIMioDqylDfIdf8gLhDGRLJLRzyOGCwSAdvMOIYH7ise
Y5ppNV1o2oOG8VPUjZpGMeBP8VSJJw6sV9L4HNQPqa0sWGXXLmDBxTb7Z3oU+653R1ChRw8ICm1f
PgwWvdXA4edD0+yD6ENIMgRYmaui4JA2dNkGX2jYadvxeQy+1sRLMigkekS/4fG6Icg2fMOHsrxo
+ZuDS+eogagDjnuM3JRbyoa7ml58B9ZOZCkIaXvzfbp9UYQgGL7bP3FoaZ++xudlzXVkWJcRnVSu
gk2xti7KzJSVcbAayJBXgUxJPPs5HIFkj9dagfHHLe8hyqkMf/2Vmp9QMrMjuGvH4Q7n7/IZ+bc2
sjwygVIWuWAgA4U447/n36uHBvLv0+uSIJcBrRFekdLahvp9cH3QgTgmm357dyQV24E3zpXiARgw
1jPv/5IA1d89v6Rop3CWU7Do0iWp+brtR5CluPa1kUs6gbjHCevia/By6FLrY3o3EsygJRlGZZHT
gslbSeya38Ns6wAB3DO4io/omBnWCxKg4gtnn0s1NIQ9gLHqI9eexHr2PssRKp+WVMwFBdb8dwPl
X+dr+dnWsiL/3/a9bvYSaRHgele1sOU0znhz3Mh9uNHXRyGrG5hHZntFGgWXwDkeW9xukULhJZU1
L+6zdmoGdX2av740KK/04MiyA7CncI91midMkJFGBx3zIYhTE6l8gXSlCl49uzoQ3bKCEz1mSuoZ
tqpJM55CMAMqw8/ep4im8QSDGac8pgulZ1LLgpFiKrtJEueuUYcHrLIeD1wiFF8JKBj+A65kS9q4
YKVFuLoGEX2WsnPOqsDPe2FwE/5VdvgqspPWr+H3gKuqCqgrNggmm8x91ZLbYJCsC88dAjNOUWCI
Cr8Xfpx95xi2vBq8ae1HG0pTxnZpotLUiPpdSlPDISgjTizEjcGXPFbKXMqNfTUsifJIv4xcgRqU
tL9LyFnnSSWbt4C6CyM5nUB0S6frK2oOHPujWjr+SjlgO6rhw5uGmSVKTv5BRWBsfi6CRU/yQ6OP
4+wpHDFyGagKoKx/BPc9h7pUJ2EpFMQ9PZUheWEfHzkFcla7sISadxz7Eo7X+jZpbXB2TQlok7ee
KKZG80nNoqKABUec1MPDYU2hbmPnsDimS5zheTl3nIklnaNVKXUzTCIRj477nPTarZsH2wBxqoPC
CeIMZM5Jdn0q8pimPtjULlouZgCnkk6I+/3/ijWApjHYKmIJEUBNDLfbodiuSb+YeULTXZLBdO36
zSdCG6gStE5VHDwgsUMgSoELY/g2bm2Zn4KJJ3Nd60mVIVAzg57hgqdMSF4qy9l0b6GK5jfl5Crb
3pl87I8D1pv344fbbV53Aq9e3fcpMxBs4VdxP0SrNjVnmohljOTUPESja7jppFjhgGeIS38FlonC
q45U2iUeD7jb/GrEQxlT3onn0LqAPesTdOw8hgWKubrPMmMBNFC+JQXuEZ90KFOHtEJi2bVeHHlg
YmBEShdIIaGqee7STfww6fvi095EJ1HVYyBGkf91P49oLg2XSBFiChTutqVI57OxRJO+mjhx1hhC
3CqCtdF0uSjAkrCIFzS2Rd9pABmyjVSFCneFMb6ZGER8Ftr+K4KZXwLlH+2nJ5gA0xuJN63sD3E1
PkAUNpkD9/LxjOp7LGR/jC/HzyhQi4nGI1g5NCWk9rbJXV+uwJ/WQXucPtajqkpKkfvXwFI7nRxH
raRD0T9ZQMXX7U+kyohmh9eOtDfgj7thhJ0s/THTS+boheT7z4Fp7re7ZjaWatDp8Bd+1lzGE5aw
tliudSyJXD1R/yK3fpJUZKCDITifnyuwsMGoU8YAuUHySzugtT5FSGrHguLCCuUsUqo/ooi/k8fb
tkCHNwVWo/byB/TSE4rPqSYpJ1DhfVZwdKmHJYJgf2DhEdZgaETSe/LrtbqCJ54CzmRf0kAn/6vy
pdrGEkeR1GvyXjVDLP2deLmHbPaEAvrMlcHgX0ydiNQ6d/MP6c8iwXPlMnHDwgaGvuLXux+eIg69
rpFIJYJLYpPlpVc3iG/a649G7jtNzOFkV1lBTx5a2XZvnn9Z5yyxkFqclMlL08RXC2jyvQoIcFLY
4SL+jhXc0oWx576Ir6+aBhcnKwz8QBc2MFebP9M5w085lh47lRJi6IGw4NQQ/ulU49bWjvOahKQH
yVsPDeId9xmowV6k9xBoOmRO0CMfM6gwLtOsJiUAJRGqqslLaKqctaUK3kh/pfc0TsFYLBcQkw+6
By2FaCvbeWgXiNg4gfCFUXVg+DFwRpAXyc7bk1lay98DK+JVP6crufC5+NxPUs9klA9w6JQjJSLy
FfuJLgVFKstUvU+XEz7PWOxhCivvTLfv85dcO1OTC6oyAAhrINlrvogIUBzvSUqD2MGQSlUU4gKD
+pBAprU2bmcEoxnXtn87vnQF+89djT1Mtao+WSunFoL3gWiU4YUFqa0IGhRKf74VvrwJy2QB2rjV
50+1zZ2p6TUl6gOjHjm5+u7LvU2S40sLAcefuAzxK+c6VkuZHwKWp1KeMWAPoGSY/QEzyihDYxAd
E53x3X6DS0qeQZvmEPP3SBXor+d/TK1TJkEVoFlN217fJ/jW+OwqguPQzEJWqo4jcGiGXf1piHvr
Lf7OdxJlhWcJVh2mWlXlWeNxHQ6zfgqbReWwIac4ZdPZrt8GgvRBrrj+x1HjQEcJ9exzh7BeXlM6
2KlQuN8vi5SlVOyT682nPb5LMhwfRkM93CDovy1t6YeItUwWHMYGzuhlQ8hkZrd7gODiahvhrXhe
i+0xlMi/RQXR0i04tkxHjc7Hl5HxU17NhCf4sbiKPluqZc9DuTOlElb4AWRP0OU1cfxCA+7FIEIN
LnUXqWzAVTpIBTqVggCJudzskSzhkDCW3WMorGkJlqWZUP8eUjw8Cn8kWgIPXW6mW3OI46zSQe2N
ITTeowK2+E6DHcDJovdrnfh6Rc6vyV2IhzqylTULyYnwYpZ2V3mCN8w/gDF+eoHTs49c0mBdAE/L
5GU5n/tFmxprkwDMlNEKTSPbRYUIdr1wCmLX4vmlJNNuWt19fFXzvJGsBM1VxQ0NNjzD/+eCL9Ec
HcwC4y7FjP7sDS0yOV2HWPoVOh8mHcdu8u/Kx3PArjThzi+Cq/chaQ3y/OFgi9GUgRwbfk+ZJh9U
uxXjZszbfFxL+tnQRyxAH9GCozTV/OIJQRRIpJB4asB4McnqJ/rnH4hzhzGoWwo9PI5SYa/De5ms
Gr5aZnxMNACZlv1PknJFRTCAJEX50YdD/brNgp1wMPsY/MkuE1+adE73Fmaasrh6Rfy2NCv0DASN
eNYQ8j/i+1qr7rvwWwfnHnFcQtWUMzb4Xu09Bq8qAhcs1hUUY6cOExKdmpEl0udoX11PcCIs6kZz
+XZC7sNkmbCK8Sutwy99FflzwaLxJ+2epxsy7i73mWWmGQvGqhYAWtP7GPFbxR76hlX4xaDsFLRw
KXehr/CL01BsbmQhiD5AKBeUpemtaXBpnjHZEyfSROmlh7bw7HQdSelLa5EPhAaSsdReP4wPCSr4
mB/kK8FNzQLop1wJ/5q5I+ZUVzSVSS45SsbilxX0ystDe8J2qWH806c8Zd5JoQ1M4gnmCP2HHH1M
MfByvedAOAXeYMwPsAgjD6NA6iY6G7MjKGnvsGIO4ocYx7I/sQROhO1NNT5+45Q4DkoqVWRrfr+A
ajq35B1C4BcYRtBzzl/2eqoy1RdNppYAiKmJUS8HQFj8Sy9p41VZPMXjeOFlTNf05x3qh3Jt0q56
7BXShD+EsczhD4mTE/p7a6o+XlddWyr7hcv7B+bJhyCZ4r8h/b6d+ijYGCRGqa8dikFBiJVrJ88t
ag9Se4KTMi8wTC/cxV9lpDNklhiWKbziDuKq6Pf1wtFcTUfGwir8ICYuaJksICNpttu1MKDL61dd
nTLK+MhmDCw0lwLiFl7l+dRDX1gf9M8/V6yB9puZo6sflJo/d6+BpAU9TT7Pl+iuMmzUIgQC98mv
Ga89J7jyDkEyrueEwxN+l0gpa9/RwoXfnGnv/jc0F/l2sOw6gAOkixbdv6cDUgoElc6VNxdC6DHW
ZguUkx+gIEpep8IuRSRcaM4OMiErwKvy9vU3GQg0kFpJfo90ffybjO3Lo/MNMyTzFnAwX+iXmQo6
viKoK8oMJHgY41WNKp8sG//RZ9zWXUd6bv7foGjGySng4wJmBQ3r0cHpdf7vPlmMQaKx9gggQ2oC
ohAUo4aNYnkKX2KSwBtScyxwnI9/B3+Z490E0PJuShCnvj4S5Lo8FrrR3JOxtDR340CvyJ9oKDFP
DAJoc7VyQP61350zGG5kH6Kwfxf7fDECsmfY96AxgOml1lhEOvnAUbw86vAR7uEabgNEbbbp5btC
N4z10czTvPzrfYmBDblzNiCuEmGAFgt6KKUKt4GLMFzJc05QwUewEv4pjyxfAv9HEhrVbpZ1f/YB
QI4Vl/9+BgF1aMz0xiQbbU8ImqepbkXG6mqhyRaGlAa7gdbkGI3rQD5oBK6SRPjeSf30763/kvHY
GuycJQ0J80Yy6MLrTlYo8SSvo5EZkTtz0tS9LPi1XBVf+Osbix9rc3FVlx5MU68xeN9jHEPiiVam
5dVyiYL44ny6bfqcDHZrxa2+lqag/vQwB/eyRoKT5KWcT6oSjQKp/oYbrjk06g4TkoK94/zAJGlJ
bAVF9Bx3nMeWLF0NpaTONYARaHWulWKjn/zIKARC5CyJxgxnPJsA6yGmkKeAO4qavp88ge+pokyg
3c7oV0fawxDXxIySYt0KO6VTB1V2WGo+1oCxSYJgxgKx/mmzAf9IKRWQPFz/DORQAvrSVN+v2Pue
YdZ3s0ZVGdk5oIiSw4x+H8i0qwHeFc6DU9MaLpeUftRR0jUhR7qIStmiklLPRbtpuW+YbibVv221
2y0wa2/gkAvhxHYShMBRidayZ3ePwwKwFUVYE7wJYjd6T+3k+1pKKVYxLSRyXtb89XN6L/w6oFrk
VtqKrTFzvcuYr06yRCGt7y5nEPwcZ7Bft3x901S3XY58LJIFh4iuWDr4pSexAVogMCdxMH1Gqt+c
mWJyjQQuSxpQnzskTvyeUKxbOda6QfGeibP2/Mh4vwwC5ErdddbDhJtZBMo+BJyghlx2jkw5O4mK
v6X3QYV9H/j5rUpJ1Vxt/XJe0jYa8oGdbsTlDnMBMZ2s2KmxPD9BseasBsBQTJ31Xa7agdWNaLsC
EU7eV6QTNYyezpxX3w4Y9CXzOG8OA7GJ/WvJw3604tQ206dWi9iLqHjNpjf9fCWKjI74Uaf2p/qa
uFTy3hXKamQJjw1zClMBkgQsnDOUjsieMq87ioVKFtljzS40bOdqPGXg5mhMWgZwvPcBMBxN3agM
Zzu5k/vKKYxATKq5+WVBgyADUkcEe4YRCF2N8zXWE9/MI3NkWMcpjg9m2FiVVnbYzdI282sINyy9
MImXOjo7XObxYlNcVyMWzbqWIrGNb6qOosnNu8JJ+5ozoC9XVmw7/Ij4hJ/voDeJZ2yt5lvkzc6I
tXxIlI7RV8S6GVxxUyX7FB6hh8SeESwaGnWlNxMW52H+4i21l29SsqtdQxtCkrWJ9Dt67cFqO/yu
6g99SIYwt1dze/AYiN6mVGPq8cx9JwyK6q5PYVHXfcaq6uXUEhY5ffv3+qVi0nP4/1LYGzREKDTW
vI6Q/RzESn1R5T43BLWUCXy4gCGuTwrG/+xLK2O51lulc9V7GA49fNufr5PrpGG+sfCm+HDpy7QO
qeBmCiqYBiKeHcwirYv/N1D+aUXCLRb87uxA7eSR+RXf+YYHa4ckmZkAjcB91RFi0Tvs5Khd+u2n
MPfY1tbpWyllsfRKOuG9gGYCluNf1YHVg8wqBCpI727GFnf/qmS26noKy4JairTadKjUUj/XKnLd
dG6EckgZBpDDgo161dEIjzZwzncmiGtKA4fDiZapB2OW0z/JhDPRoZ/+lBQWFuqzWjEe9XioUoXG
GHY7YIOV80K0zwJhfsv9dBr9+jV0A9cYVz/uE3Dvm3j9FUaYQNIS4ZClyW7ApqGaULbtThR9Map8
6Sx6OU/GdCZPdf2EKcZbp75ivSwgPQmIyU9s5PbeOJTlQD0s0NGqeyuUxF6puzAZzaIhkK0wwaeu
ERayNhDQtzrHxIIf2cBGmFVqcalP/WGJ4+/RJbwyF6SbGRmU/i1QgumNWNC5Uf7nvWCXGwT3g9I/
3wmyVG3flXRARt/F0QwLwf9CIfPkiqZcV7mTAdxy6DUSbu0ADgTvkPGttQWOMm5LQU36C93hcAcA
ww3O7wqomxVVKePhh0KD1bCo6HPE63hy4woAwO1PqYNdfFlF2MH+PyJEQ3T888SJU3hfka0kSZiu
I3eMJGkfJNJBHPyNrf9MItgC7LZQaRESNm7rDxbda7e/fpEDT+7GcpLOEoBE7AtiX+j/swoAvFgI
0dukTKdKItAGLX/rUlC69Fjc2uX7/85vZP/J27/GsgcurcMBOVmh35g/UCCK3lbQsL0NQH+ZHmu6
/K2StabeBaI0Tyxdqx/6+d7ce0jzuzyXWbLAmnatuRy5V8ZDy2NsUnSC59bQCM4lmksoPinNV7Ue
6ZMYTZwZ64+Yr4oxbPE15IBLToXImo0P5Yvpl3O3jpIRTNN9RkVKDxbP24wtNEzN/xQ732WF9Z7o
qgjxQUBW2NrnDrEwnlX1cQtb7Z6QgRLD6+kka2phNWBhL3FhARgH+hCq4tEa2bGokHuMIihTQsOE
PTukBC/YUHuEFuYsnm/URawLOFz1tndxCTb+SduJegjMqhR4ojLmQHwr5Mwcb1UiYvqGGq6EJp4I
e7iwhhnoOSOi1KunjA1MtkPzJ3WtfTwDGuXLEUUDU+dM9Hq1LzJalI1XuRvJ3N/fbeVOPsjgKPxD
agXidlcYcvGwP/i/jt3Iigd2iTgomD16xi/DfYBZQhxOUdCe9RkzZKkIJ7TFzPSyb0ZWlOrqHlW9
tatuo7awlRjhAtXPK0RhVx8bxBbk1kLGuvmJpEI+RJxi4eV9t5D/ZzBrMU7cIjBnM3SIP4h3TTLD
G+/MMjEe7LufXYvm38V+fhazKf5Puh+6xunw3D6j4ZCTC5wJqo7EUSc8GQL/j6yREuE3oIvxmEV8
ShLJ0O+BF0eAeNtMKlZOCJABTv8G4MnxWQYmcCl9OgvLyLp/ubUnbQBUhQxu4qljGUvkKurbJ+YC
L9pb8JK0TbH+xMAuJE7EyUYE7IJF6ottHuOmZZPtjwHqbFUNAMDb36ICBn3VZG8wU1SsY9dGy4/0
kRZAS8Xy4kVtGxSRUmnSvhue+iTbD7hLn0/gp4nazLrR87+LVfxd/ppu3bUQKuiKvp//mClXUguF
skxsfWYyArwj3RtU6aUA5CDVxx7MPaqw+LhQZ1DUc9IY59cFcsD9WH8NLsYqnYIz0EAbbeIrgMqY
Ns3V2zXLUlMtpEGdqzbjqPDABAsTLRvx68Lt2f258Ln+WB4z3tMbU+/dvPZAo3PmIu1CCfpGIvy7
tIsN5y+Tq21EfrFHvmNK+nIUR8QQdQgo/WF+7Z+8ps2NqXtdX8rjjzce7nX+2JslFHdqROXaDiyL
gZVTfysWZa+noswvh7foBuXEGdI9QL6XeOyLMqDDOhitOAn7T5W+iHDF1CsUJx4xGFfxyXqeDJB5
afO0qivfwViGQg5nukRQPlx1WCMHfCexQKJ+P4Q0tddNzremOyqJparr6h9rmYIT6WwIxlhqxbyc
kE4KEMYZzQ8u9GRQavs1uSPIMMVZYuJENk2DF8gK5U1tppan6xN5VVbqFooqMpawql1ZrK6LUM1t
9e+M8fDSTignJgJzUupp6KUD+KEVlVpTJicoL8g51okTeN+Szxw7Y9RZgqXy4432VktJgks5LN2l
Dc5srN0Oxubz6SSKWXzHY0wTfLFlJjbaVjxSzQRWcLSApdNENAQYnI5bsxTeNhiiPu20MQq/R6ex
Sjy9WpdJxv0uQI41lmjToWMye3tY1w2ZCTm6zLZBdiOfd94Soi+jFlgEhsgKWOtrSXQZp5x0TMAi
ViCVaupyHU6ETTSwuSgZmATvZbg36QCVZ+hPNqazgAh8Mi+1oFqKj/LmWeqwydGJplBb4DEiTq2C
31YQBMQs5ZH5CSGGwjXBENLB0H5ouHYjxSrHjd+nt4cbO/DhDJx46p2QQ3Oa8Kjwqa9zNgA8kEU0
VTmFSSx15DC6cLirXUWQDa+rdHN9lud4sPfSFXqgKVkXkXwE+e3XoF3G51J4R0XG3qcJe/rAvKGp
aisqGRd2LhE3XUrK95Wm+zBAgKRm8fHHTUdjJZeSZ6C3YLQcjbPb4GJ9QhI2IELxh0YghWw6Nrtc
BVbM1wSzTVMKw9kxMWi+drsvO38hHygem/KTQtEpEZ98lDZe04E465I3FQ7p0N7YrIBNff0TWJns
s0bu+j16f0PzzQfckkz8CUl3W8vZsR6z3ZUnJAwxTJ0BU2vAfJ9HCnjXl+zu9M1eJR5MIRBsuARt
axPmVlpqbZvsCQ8QLSeC4XZ/LHr6+3Z7K5iZxdTxDTniW2Ezhb7AanIZ3+sOhk3Q/Oe+v4jIXKa1
LIbh/R8P71YwoP2jN7w5wooommZ6snnYV7Uf/+9T7NFoTH6K0nndSPXvpeH9tdYWz/6dLkw4jkrr
qiJNo28Ilut0rlNDjyi7rpAyBZWf/bHnf05Ovwv7dueKSxmg/Y/1pVS99enK46WQggypDmzqZj29
nWfQMyJVF/4uls5w6tF+ElLSclYnipjc5mLSRbyumRmHMqsY94OBTyHfwu7czm+fc5cDiP7+wAXm
X6dB6sBNYp2o8cPXD1vrxDhw4endPGpw8Txnd2d7knKuv5Vst/SJKsFZR5rJBm2CSJ+0sc7sWyt8
0DgHtKhu50gWp6nTzUGToWfTCppactvjJrPJD5/ltNn/kuRJ26R31mGnFFV+I6KWbtPcz+A3lseh
4jQ+ttNo2jXxBUiPcLfVK8vY69QyaOxbAaWCG7LuvX3t5rGe/HvjqMAK8NJZ6AZGSM5/pSWDQ0mk
2lKfAHDiIB5r141ootMnhWFwVZ17i4mcdK0r/bdyV/SbaF72VVthSnCWVB1bMGrVcfexNPKcNgAm
vnSiYnoahE0VHzj0KqFe4X98d0vlbHwt441h4fLD+6VgDJY4+2hPYwpzyGMZVzNvrvku5v57dg+C
YgXJkchDUpryaKw3Jbv7t2JitzMqqDqMQcZ4gXrBy+N8V8JwMrIlzeztqFDKTvhQIQB2mxTZiA61
cc8rOylvi39xB8BP9sakqYScxqMpwkTNbouNGfZkO5zm5nEXyZxr52dMaRQfPdDSTYaI4nNgri5L
fETiYKbl1h9M0Q2CMRSR6pt1BvCbNEROSiOAgXMApzytjasrz8FRmkGYWGHvGhuAIpmmWxztZSXc
lXULna56FnZkSAb55v/XhsbHl1UqbGtG7HxIH8vIu1nbEgNbY/FR/aL4pDahKVpBiyUtR+4RoCvF
MAZ5iM9eyi+6hgnYMV94r3DCMKY7SPWvuyrj7KQVLmQlAzhr1fvb9GjnOrLJLIBdzGGAYp69ZkEU
hMeV47Wntx5KzZwhhkCuuDhSXjHy5O2/IRghrTdfB/gZSXExVdH8r/htmoE5dq34PMLnX+R8BaOR
7z2y8DplIi+oIZafP6njBIUk6ag5fWdgK8Qcnt8VtUdyeVbCq8kMnpk4TnxSVFS7k5I81T4OpVAz
E9Y7dTNdNq05I/hsMCjmEB9gUiMKlxFo1CrwXCq+9erZ0meTGe+ciRpmm/+AVWcImce8/JiLlYeo
r5TXZHEwybJ9xoNRA7+NALoBDiJz7KYE1vdni9dlVEVPqQeM45U3TnTCLfs6OaWtc94dQwtfWUrX
YONK4qBAbWZk9Eo8CBryWdKR9ApPOr+OagKXL24d6tX70x1keTjxgLa+T0EN9+xNX9L0nGJljWNo
mFRvA0uA5A/1f7A/5nmxeyvPgwQSAeBVyf6teFFdM6JkZSbeU3MrSDK3a0LmxxccP09hytDYHNBv
UfZ17IQQs2jm18T4WmGP+s/M2fzY67PzLLQGk/sie1uREKkVBiXpAwOtHPmmTEUzSsO2zHcHpPTV
4vIgtixp587TCGpyC3imlUxdCAcHItfbMuw/2A0eaIK/h0WDCl4WOMkqL+49zCEWUCj06V+YQ10m
3VmZ9uzQ3FWMbfwxj9lFaS18U2mDY4CMQLoZm2OYFPSpHa1nXPP0y3rJA47/HreJd/76qsYE1dT1
tl0OC2mFEKvDaJz5hZl8NNpZryLlkODwdNFLnT3GYFVkYx4E0rnhl3DMPLgB4iPg89mkQ/+6FgIh
JVE4nCrsk4RNDKrfG7Uq6vzwP0ABxD+3BvmEjZxMRtJkkSc8NuvjSsxR3Ldbo2v5jYmnh0KgodEL
ciRt4MCmfMdesfKwBKg681tYqgeHlawyyaBOc01vEiNsAVPM3O1S5LxxSqgVAeNMf4Q+2dCprFdB
gvZA+VWuI7tRbIEmtGvpL9GV0uGOdyMYvYz9OPsKiJoO3uwnBVwb/2WPPtMb71IZyfliNDRqQ75x
oLXvXNuRqcUfqPSJDl198r0NiAdolf/Ba/ekAHYMM28f7M5hQtKULHSz1moJef27qmy/xkkHqhhQ
hvMfmyiE9gcYel4hgmV9YpSx6b5JSD1OhdDFKlPcOY4nhSiYbN7fSrYmKtoSNPGeIViucWA6qzxl
CDElQ1f/D1Y3uQMO8Zoi/UhL2BZChBjoco0hXoKz6cQPkrZAeo+dgDKl2R2uiyaiCbULjkqBiPte
jJlzXa4Wx0LJYBdpOCCat175nKphEvhnBGcS4to5ZWzj+JvHsCXiakNY2x62ng68sSbCQr4J2Ua3
CJNX19frdWM0u8qyP8sWklPjDqyAQnJm1a1n/9jxcNa11ke7v9jrBhH7ojnddWaXM2GGrqmqE/qt
trLRSE2kEse/IkfrvDNnbJTKOw0Ngzc8RhfOjlIvsaJ5Z8S68lqNalUvMIt4mFEJnA0jphnu55Mx
dn2wwmkhsJVAeMjKuAw8x6vg+Tg0S93rcqBZVsizxNdpBcRi1O6gqAGf+o2sgZEqzSRVdUJYl7GD
7FqSJv65UWFcLDPVkbrty/ShzWpkcG++cx8qUECF/5j3Iy7h3MgPepDwfkZ+soQMYpXQNOUbhXSu
ULbfCkGHUEeExGZ9ZshIlm4xkMRw4c+FRjgxSXdio7ALnidS3yLcKwopm48CjDwV6+NXdjdIRmwQ
VSVbbfkGyyzl8vnJ3MrcI32c5NXY/rxW13aCl1oYrY4NErNSaQFKMhI8K8f71LizuBeUbMRKN48r
jZsSSQ8drBS+DLQOGd5nS6KAKS5k+Jij1HoJSplnPUtrqsmIsZezPt3P5f5QwkAL0nuczj04lsxb
xhyKFymJube3tEcd75yWtYP8nCh7bQVIy9nZEb0TR4US7dLhsqcZEIzpKLXSJMHrQQyU9xwR/hvA
SJBWQVjp8zdw1ZjWtzT6WjBiwuBJKJAVBFRWoYr9G87RTP7tJkOyJFgQ7+L2soopfJXFELh4LXfK
95C8/UPvk6tlZjA+IxjTv6hXlPKJsG37hHuFMOIlDMaRPRt4asfnBKY24W9OhaOwp+awQO+a+BFy
0uquBd602anwQ6Xk2lzK5sZesaSHnIk4JaCN/3Ylu9quOJ/jhE+Cvpli1035/2GOT7aYY8ZP1/ri
RG1/enL+J2EP5PIUfjgP2z0kianV+HhRvzGhiAo0uhMkT2sbMMlFOqwNIio171Vo20M8nd/4uvc+
V1VUCtWnriPJUNk7cQKxeKbn6+OeAZ9dS+XNSQP6UiUbn/q9rECJAWhmbBj/FBAFLiCcjfY6j6pj
3hCs7CexVg6i2mw1AgLQ2NNKK3V0dHsIqJ+4Q299pMXRPGHhm5T+RZEC8rc/JcsyrG33NrB4OccN
5jqfFMgJQUjn1dFFFWAnLAzh38DMRnfgbR04jp4X0QTahyEuPd/+Kkk1jRepnWEZZwRBeZfe4Z12
0JMLe5h9833iBOs9FtKEvobMNbN6zFuNjGtstT6wxBZ6O9XFAKsHLjMV76iTEc+aOJ/KOnFnjEB2
m9533bRWTizsYxiZ7rrS08SYz/IC8ZjKbJkEBbqe7CZDd6L9RYfjWVbL/DNpDtlErnSB04QNH64+
5Py/hZ2bvUFFQHAQKVPSRUws+OhFQF8DDMU4eMSWHYIO+Mbm4+PrldR6jA3KynuOKu3XxwxBif8g
4qz6sFvlIufg42r69w5PW8ZVAgkzF22r6Mq6EMofvLjUStpLjeROKtwdlEE6Kc2ZRjM94iXkKYBh
goV1qkWwwQBzPrI5GSz5Hk7ZzUNEHBo0R/6riYHqMhl/ycsyrHf8ENo7TxJ60vbGpSs3bXXTIt2a
g9ptupitCLc/4w0GUvVvWYALUTHIVzx+61xyNn0iQinrc21f13aGznDgR6FgzvWelStXGU1/oJA2
rQJZiYUP+pTDNdkhufFGxUAnmgP9GrCaOZpTBxa1r4BRz7XDyD/BTu30ImHlKoioGqiRcCUz7WAq
wglxKeVa8sWeUg++VaIOEVQs4tPyy2JAKOlmWzQV3iqpOmbi0kJpoAW0Y6jk1htXoTey8aTYB+8J
CJyfnzP24gGDvbZC2SIX/Q25LNjg1D8JFOEMgKh3yw0qJ6WmhwJjUNhXAlT4gCaOOExc9mvHOb4+
kFyTPJDRMdh++r+jP2wZkknbmyDK1xetpHabX7JwfORSN9wv46+PXdeUOlRk/6RFpUl512vru3bm
4Oy3oR196vJYvvR7S3NtvPn4EzINvP/sJJikVCnKFuI1TVEFnfTQrZxpf8EzPWwBmw5X7AfgZmyN
bvozsIwUEqDku9GKaSezFVtKt9CA+/adukgJ8h9e6xBxpJbWxelVFC5SphdHjbKMpMdKwRGZ3d9K
Fx5W+dpBF7Yx8f9X7VQH+NDZ72/q/SH4PtzlaPDcmM2VuegMDGTuVTO8azHTVpvZ3kmaTyJIarOt
ho3gB4FUG/U1F+0RyP1AlHkr9yvlpZ9jpuw85KFf1pkhKFHmXrMJTmmgVD16xG4nnckhzBA6pOew
uAgauBQaz4OzYzmC42qqwXQSEC8DZ+d/mfRqE0y/oUAewwuHmCuM7Emz7iYvc+cxuQLWAIxIK+oj
1tK9snho9IEN9LpooyuaJAjjabxDCdAD4ZGW+OXdBSuQSkSjnTG+Ap5eit4S7oULvO+RUU/sI+Xr
h/CJkoO1Rttj67Z95BrNjeMhHhP7I7EoiA8ugTR0FRILU7cgLVqEo/j+sYs0srfovaKi+zXs/c77
r4eFKOOMqHYfKEqGNi1JbEWy1aKP0orFEHgKbZuBOITZBw+4ML+Sps71zy8KUiNF6emccZ7PR84z
sgeKsp4sX37GylVDmDeMWvsKDVErQL91x001lJYkb+nJFCdb1CCkWKmTgJFVhvbkWU8LAINKdWOC
7W7y42piDtMC3dKW9/q8IkwNoq6EgFh0ND/F8Drunaco5Gl6Lh6xpJIGtaA5SmXLKvxjvWQimEee
idRBAMkio2jx9HoR82UAjxpuILW5UfaeMS1pBTMaUmrCRgfEjyCoBWJrHOnq371PEAc7m99+sM5R
qeKLwmQQe8KAurdYGMezpAg4tUmD8jqT0bbKVd4H8YpHbpqJ85p8c5VWJelqI03PgrEH7C18nysU
/R4Mugqq8WN0vlOqJLKzsmj4PvkPJMC1wsHRxrBRytKsWs6XEesPalXr/cM1kpJB8RQZRkeOh2xN
uYhPgh05zE4/DvH10XuaLuHudyA2/Yu49al3YVUIam0ByIxrhxwuspug1el6e2da6RFI0ZUnN2+P
UOgksxYBMT+4WdHXqswO2or94RcAqHsv4vuTvDlRYOdJx+ml7oeAuofcahkc/ezZIru4HZ+J+Noy
zYS6ccznwXjNHX3Us4Gj66iUlg+rRlRauzEZBQThmwVMffPEzMPwW/LCT43im+SGMXVkSMlBbI37
F3V/T2i1Pz/LU6ThY2Q+W4r0LYeJP0cDxwiNQOv8xxHIQUHMYpXz0D2ghEc3PVtM3kO2b0XdFNQs
KrHCxviQyUtu+81Ug3cx4npxVndwPfOM1s1TTeiEEXj12ReEssxQxTkQamKSn6Vi8VexRwVjGn/h
vpuXN0A3AvNdQW42s1XSk/YSrj2MPhuOH6xtcFLyBkP+KSjymgrySrIAyBaN62mhMeHM3AP3+hiD
iL+P3kNjX7UCaiFnrwORO5tukxbI+AW4isEbqqHTFtQdPrN/q3NC0k5ilC5rgy25VpJkSuN1lRt5
cKoUelqMEUGuBbqp/txGH6M7lW28DUymxads6SIaQ+nqdChNT3frZVzOmAWXGrjfhhSNl6LJdSVs
GtS35MP8Jzrm7X0BiYzVd8ENlqXq59Ep89DpRtPtBUfFDmi9IDuPo/jy2g9NasDXV3JX8+Ow2dXy
9NUn5+CUMyZrYfEjWF1trAJaVjCSioGEiv5aHUjuhtqihi2LNNDGehaNxuhyjjAF2YU36cS/oLCy
nnjFCtRgfFUGTTtUuHtnvYXxBLEbMa/6usxlZvjneEM810INHCiVf9OZC6KF6Bqie5hn3HYyOOgp
9hKTC343Awj84TNyXFt4gU+tXPXw/ZiwI5chdu+mS2m4IzDTppMQi4aBbIGAOC/M+vaqzBZlFkwG
wS1lBNPjgEnOc7QquC4cI5Oihf82DxrewyIRtzQFT3uaGMbnxALhqTQXJic4aKMyl/wmOPLi5vmv
yBWpFk4W0m4jMdFCBgGTxQJAjs7Et3CmGIY3muu/x5QLsGNMoEjmzbxq9PvrxJxnR1SojKYv9BFm
oR+++QeBMTbQPWzPpDx/5mEJbzlLATuCe5dQq5u9zJYmLmgoblxAFEF4+mDZM73H5w9N2K4v8EJ8
Uc+8MSmTqM5UJD3FgZgIUqchzY02KX2p0ieiRjJkRKGpvUdlkr4NloqH+UL5m1dMjFZ4xkyBC0Mv
nOQ6J9Saht9cEvVexYxqiW7cYLcqBEkkeCPGTMeFCtFWZeXd3P6u1nHYWc2uYJ1sw3dpxtWZf2k4
1glINX5Aii99SoIJJ5346DXLgJ/F/aShuAQa52vJKFyr1NSUiB/YvejJtp1EoS6xxoBz2GpBGK7r
FG5k4TtxCaUUQDVhOz4nAHMKR4CAmDGIT19XLSM4fPRX0Dzo08jwIk3rPQJoRlwaawcM99yIjHws
q9TJcsfLN2Ozvx+9UL4qehhK92/kzwkGnlY8H/X2IsumDt1VWMaQ1FPefibL7jM6fhXC7ysWQaeO
uSLT6LG3NIpEhW7wTiS//Sg1QrLsJf5aYmE9+4gkIsfyTn6OgQLLprPhMxFCM++Aw2RnXSt1xzYf
tc64KTcEvEPRIj75TmiHQGPjr2B8Ebm/t1PvrTgzNTi4vXXtwhxOMQERIu/KQ57WxGcgEi82Ew6k
3GWavjb2SA59hfBLHTkH8oNGXsTS8YdT6ZS8eWBJm0v/MY0drHZb0c1Pbr7Ecj7ZEchzZkgPSA7u
VTzaf0CJuFxCQYSvnDbOBXSq2VWxR1qUbV+mkZtvIQ2OMdiaw8oeC2nXK7jjmHJPUwpu3qeM78kq
Lag4g4l/BAblJGHZXDTjYuyVHxgXDb6SoEZc9QbRUhAfBOjOfdbvHk7HwXHwh1BdLrMt7kMx+SxV
+RxvD1gRESnhUDWDMyZlhOLzpc1rVsEJcbmZx7ZfvQyKys80NzjP2472rp5l3L+JNCHozxBZEs0J
PcA+06wY8+WmSXO9KXurmxATdtcqLMRuXeshLf+P1WkHM7xYmAU/DFim/Rh5ObP1U80e3ZnxYOmn
d9iBIAetFSYA1wSzSn7laxHQb8xV8UKQEKvjz4SuSzxatFdpZrd13RRnlTPrxfQB+RU3v7muLMNd
bUtAMwwZOmfbPAznvumJK0oFuuSdGnnaT8OB00sWs/7a0O8qoHe7EkD92VEemFBOJBXT6toMDZ2+
KSSpXVOSYTopK3eMxrlrjgk0B/sHZE8UDVjS3BvzeHshCDB4wLiFzv9tAdz8jkhst00C1GYpCBlS
lRKiCPb36iu+JJpoZNjXRomwu2zfl0vkX1EIto+lYS2TbZVlGAzyAN8ofDzp6ot4/zBA0unjoZon
zbisrt4RkzdfRF5vB43A2l22csX2fR7bKTweQQbQ2Rmp/KyNH2vH+OL6l4qt4qsMc/VdfV3qrvvk
qioRlcGXiW1QRAC/nhSv0nFE66cKW+gYN/IlkXGsoB95VwLvOZuLzKxWmvrfCBt+zn6+pdD3QSNp
9QNBbw5JAGblFPdvVZ8vqaITY9GidAnLbB2Lm/ZzFvVW9FJl18t5Mj74l1TK+bqZ/bJCxygjyE6c
5nrOXDH+/BJ6iib4s/Uyi1+QLzfksg3UWqzWK85M6AYbpOcVqjFeJymG/a+sFoPgH/DQOko2mYUE
JT8TiIxuzZXOzUwFvKB3zDZal5hMwhPy3ruOYBYhPPJiu+uqshvP/aubNJ8dKn0+sMWhrIIaE9FB
jLf9CG9NOssZxZtFcBm0ZnvrxFueNmm89DXbfCqjNfakRH7QewqlWnL8TYiEC5cEB2BrHL0eoxmP
xeT+d+CWK8jG9sISA8Esmm5wyASg3hRI4vVigf5+EUM9QIBRy5UTGLwzgboGS6TGki8Pl2ldCqZt
BeYz6vda6tEBHhdMovRgVsdp/QHXaxRSudbgxmteIL04GAxa7o5rMStb6U7qYf6mW15co3T3cNu/
5gFhUu+G/s7PY61pUNra5QlstPbIdFh8YJ3+o4KxcbHGYacij0uM6q2UAkFzDaNOtf/bBndOsEY9
j+5+LaHeERIDwzdtzc7rDK5juAhp5xLaW3oEhP5IidRbCBc/0+70l3mfZKBqIP3aU7hQ/cz7+WLj
sQo5+nne1iUetYKcI4qmYn+yeaZM5myYeSGyjFGi2H/YUh4Pbm+7UihIWSjySgz5EuZSxHrN23Ze
5ugjFHvSIvwzc79y9m4e22FUfw3jkil/5+MSSg87eC0FcTMTYdc7Ohc4xBXEAmBfbUpXUyKe7fPw
02jMZ3OCnidFlmylwx68PkLWwZjFO0UsCE9Eqcsb8L+Z9uXhTZA9bQRWFs5c2gIcgJIQd3YKSbkh
UYbtNQ5fT60q1p/ThPpMRZCCU0gW4pJ46hjVhFl01GK6pW3LUKe7PLW939BLdZLxI6bQT3CH1Ui7
yfWUJPUlB7wo0QX0odCUHdj3tdU8VDYOAl9DM/UlcZHblUjxYzUu4oX5Fo/C1vTfauXrngiagf3t
j4mLexOEjD0KvUzw59wTou5DP6Yqu4qOY1EPSBzOdr8zBdGoCCbZRvfzfC9/4pI4alEObe1Wgs/o
kCTeB+DYnHHiBs5R7ZeAXqth9KEGYXJAnP4PKxPHCjKw1YWtw/ZTQ0XRdltkCbpSzLXkHgY34yxw
PaZ/9OQM2U5VhDbpxvbFOzjOZyQd9XJMUeOOT4cSKmtGcyrpQGfDyDW9kEnWw4zcCEv+IZFNiNqV
LfIBoL00c0b9xdz5uo45fRyyVDWRYUpOnf+2TScjGxPgW2g8OjtZTQHlY0qn0CsJ08wN/LOnRKtU
RpanMOt01KmdgNfWniEvN2yOvAy9yvRn1fQo5HK/NqHsX9qgWWI4HwjdAxH3Y9Qu2meBXv+uEVhH
bpnv38KHSjJgvu9QpdUYToBoXYvy1ltMwRB9Ff9dT+8DDmoO/mPUZWrx56IZnomuemJ80dweTle2
7i/W5xTH5IZsG04+f4y72narzfTuIEgQGbfimdAT7WEhKAop/gQJOFrJvajAPjsQ20tLF9H4+NzB
bmXqJEnvVIK2MijXwsHQTpd9muCFBrxmM3pZ2Xt5uFoytWjd1OLduefnQd9q6sGxCnC0FglocTK/
Zes0+FapnocgMMvQ3oo3kW3kLNbbHE/pEB03cT4KUpeleekrYlJjoBjJSVrA1LjuCyVagIrUhbqQ
On+RO/ky1gBBqvLbhH1izDak3fsxl4adhAqgDJjHKJtQXnDJ6S4MRboRX/K9bYA59RAvlGDKGXEU
ml+xVDnJnWd96neGyjboYDOp1K/m2hJ6z2PtjAWImYBoNn2e3lFDkdCr6iBxyYDkFx+z57HTFv3V
ODJOvzdPuS8cH+KeuxnEXtxzU0bgBtQ/1WxWCnsfN61ZZxtL5nWFIEmeaqdh5bBA/8Uxqz+deRPO
rpl5BPrmdGQtWcnR1w9uZT3LpRYxcUSUZ2s6V3MbPe4dQsrJZ2Vc3nkoJYMyBoba32LI5RteWeYB
nshfkjJHVtKc+8m+XTugmz6gS30nUYlgsYQKV7ooe31Le5hw+J54GAefPg3oITtamMA2mILw8Lcx
mlS/ZaUNtz8vbvl7sS0Ttyh7n41iHlM25aLMSI5dA6sPHp6DFn1EwAbpnlNHWy+AJWGJZ8YLoUKY
rm0w3AFnkSaswsTqdylIN4NV3A1DOd/JwLn/v54wRe7IjogWk4/8xbfMeEJykLMdsU/Bpok0h5cp
QTvwOmDU+fBTIJkMLdnZV2xg5n5HSQegJ5Eo2IT0As/lz1e+7SMcqnT/y9zmbzc46TJDKeB89Fpo
HZiT/5r4ItUFogROJaaxDvVF+Oj+aVLhetGJP8VHsC+6ks/nJSpaYKyrKdAUuDrUGNFgc2ORHLd3
oQTd65Dz1ThRROAZLjy7T45PYXayda9V9kr6X41Frx4ZfhQBfudiQ+GjU7ZuRDO5YrNXWJld9kZB
fk6LuBAQF0wxo3nmffRRuuzU9FYL6G5odR7sNckCGo+5q7ulvuojPhy4wKzW5SuKXNZSckJz6tZm
GExHQ3LOcRg55u1wdZlrAGCKOjdiotuEm1iIJ8speJNhk45ssi2A3qe65h3u3A4+b1LJRAre2f41
Z9Z3XjpYtxumHrKPROEUfWU6KfoOjR06LjOIc7q02Pr1bV9qHwk3pW3ksJgY0j/YF3lW/2I5+XXz
EwwmpHRDeeevAeLg/TyA0+PSQk2TftJT49io3biY/K2vgArej9uwUgMBj0+bLmYdjMT77SsBcH5W
kVQsxxlbfltEVYrOkBzmxY+6BaL2VkApswoEA8dFeJ32GaP5mqTofhlXq1KWJc6uPjHF8bDn/0PL
Y826aslTjNHOijmff7RHfwuXG+wS2U9a8cEhMCylTrc7m95R01+SA5J32bJph3mtmkRExuZiXSpl
HFMAXMupjQekf0xYTdfHJ105nZNInXPQ5WYS0lQfhraWnOzJOEsPjQSzvz5wRGrSK6XA/flHbZ24
HXnKxeddjWyxcPjZ5+pk2PAQrtbDvao6qp86nYdJGMRFZsnd4pgCapOkcENmqqaALdZB5gbravO4
T8LJh/JTWcdoho8s2FfWo2HExPlG5jNqeB6PVJWsMQIRfFt1MVmiL7xkSRrk/XcfsjoxPy/tFHQJ
F58SASmEVX51k1FWnJYA3k2Jz1u33zitMNXt/FDCRGrVH71cwBtcNsznRaBTxwHnnpvOqo9MppAN
IKhwbwPwPJI2LTVDM55QcEnfptOx16MJhhhkypswDkEpXZu0UfXAP/MEImgNaTiCMFRyKKXEiuw2
eWS72YgdmM0+gl413fenIQS0nlJ62+Zy0VX21kwTPV6ifiXX3nR+Qu1du4u+/3jXEjq0dK7WBXxH
CUFaiWNUhAlfYRNnU0tdnXue/ANn3Qgu7/jzGaiHfHZFVBR7H5ht0tbcq2NhkcYA3eIOErKZMoCx
aPwu81w5R4NAXG7BMy2Um30GVyVLhgg2xOGtoZzj9AHN7vGAa5/uu8zhcYew0in1adHowyD9Ox4W
OPTpecfRMoOrCl2US2wPN19mLJ91sMwsyNrpdC+JfwDscsK7cq/R4XIKsI8C1HJrYxBMtCbuzW0m
cNK29db8Na8E9q0LUda/HxQPLUR9Sa5cVdFsua5rBOpA6w9og1UUIAEjahSMND6rBa278qdQvbJn
AwPp/FGzreP+etbca8DgMqnf6wvNHCdrhzXjqHcMvCu9yOUbsbn5XVkX2BjGhpqFWFUpCLreOYYi
TxkFV+hrE1jYlrXIh16OESrnItwAaSiIIgjKcgGmnCDmzKok4WHDDwD0nahvt+p3sO9TqHpRNG3M
K3o24JBi5ZJ3ag6a987oiOe55rr+NX9DgKdJdnKnE+YAanscZdhkxwG1U5afuIzePL2f028UExUi
orFbWWDsg2yptv8xthFtaGiFt2pC61o+GQMJ6SFYDPW3okYBWOALe5TgZWCcxCrwc3hK4joBjqtX
4hIGQnA4AsUwwCmXA/C6lv2ME5+UDNdth8G6TyQ6YBlm4dyuh+Y1k2n4ID/adNQ6++Ttpwcrwsso
/WIp7qrDE56AFrtr8jft+90qrORKhqDhyepwfFlkE6hyZqA2oZEY+l6JgTlmt34qkwajXamVnss+
u77mr1TFsR9tQZb1tb2WrT6GUpVl7Wvk/SoQzhcsZAzAA/as26vUDhB6+MLCvXw5vHdyV7SWgcIM
H9CWqJ7eL9dTgaztsXExdLZQZJr8iEJ0p31Nb/Y3ufkcNnmJWgby8o34+dsvJzRRPMsw1Zmhku34
2SXPlb0NknT9dE/9ctHfIXhGLtlxzxJ9Wxjw7haQLYsvdZCoiJAZk6yw04V6VGY+EfvR0veBZSL4
F5rYMHsW4hk2H6xP397SmmdLig/qjgUn2QaLxvwrDtDiOlyDq3AWJzGA0rlG4SvfFdekQzf2w76K
Rv1+h40okgIc60uHH0anDuCbyJXlJrre16wB5Zp3vusRZr/rFJ5k6s8x4w7vcLpxGqtcvp1MNqwJ
0oo5bbw0oBihZ8yLCOrwCzlLHuDtx4a4lFpepzQBWeOyirGhf/bd6VfBSD2tN6AIxTvSRPppUyDP
fR0gU6X61aH0kG74JIPallKxjrkU0NaLla5hHfFnzxjZMCcXgXmyJC9/5eHr6/JLFH04FA+4+9Kg
J+DYF2nnzUtO+SN04cJMJjzJsPd877DYxegLlOWY5ygq6UNZOtKnagN3xqQT6aLoqTLeUMhjBBNG
NHmpSQNwTmM3MT6YsPE4RocKBB7QQaldwiaWpPCjuayg3MpzzuqKzWpYkawX1AG5FSvO76OpcTb/
RlQiDZ3MFGlUrjwm/1WjOdxfD1zxYD9U+iR8iBnbFA0N286eYPU/K6Ux6TdpExjHwBuhLBuse4zS
WMqF7UZVVshl8On9YZbVZxLUAoDaY9s8/PisTQrtafJNvqDbRWAcwVXpe7O/yW1dbv8UomqhkffM
VfDnc4hp1hlCwoqxPMUFWz//mMpqkVJFay45Bd+kIyV8XX5xdfnMOtr8KYCRnJijS8G9MBskxcMX
4dfMhPumTX+Lljp745FNlMrcJ3viIFeMfaJYfQrVuaY+yU56ijJ9v7Z0xdZfJubsuFkZ2+CpZ+3H
vlV65PjvN27mNC0Qta8CAMF0YeUO312aeFXiy+zczEsxnoULOhN6lO9QJk0zMs0E05AC/0s6pQZB
uBqu/ClX4quO9Kw6a/it02pVwJ8OAEYPojpSD/Tkh6N4C3Y0VLcAvq0QfBUqPl74AqOCiHmfrJej
vSFLvpZU0IhU9uBRR3JyUiB72hLvSoVOujIfqy7Wj82QX62vE5hiT+qNSznR6SoHqOD+/wlEbHRB
qTjH85OyB25rIiIL5IGHptjW3X4zxtmAcdNv8nZP+5d+sdzzgZcGXcpy6PPk5HKf3GCb3WldPwTw
TOVNlk+NFl7xDhHUWP5SuhUQmb1UOLFBkVG6Lx3MIg+MaOi7xOqa9hL7GkVlZ9ia3izq7t1G5liH
66pFp5PdkaZ0/NZlhTQIdCJA/Er1MRIRQQWhgr1LdkDnOQghtXW/7rU3PhXUC6kWlCntvQKOz9iM
rNe3fu0Gj+ApiszPO5mbMAMy/U99ZynWrixdTAPnZWRu//yvolumDeCB2/9G9xV9GCszw4VQ6It5
t8cXYcrwU3QAKEWmd8FJapD8ooiA7ObfDuU+uGX8SsgPyHk7quoVTEzNmKdlSfXyHIymqeTjEVCD
V52n9CJHhEtNSTZX8CLeEFFI4jcECKnrBYuFI245+kFRPIAr+iTsyIZ3EL+MJPz2UWZgpb2pfYKs
l1e1TqF22xPXgMC+xKg3chXel37Q3n34vgvuB872XVkKr76vwpMJvUsGqa9wCei8imWkZ6I8zopC
h2mb/Q/YlUKmg8VBfsu8VungtmDKjwTrgjxOketPWUn9AYvMHhRWijxeQH1t28nOZgMAO0xpe+Jc
w3U32VY9wRh2j6WrPr8byIFtFT2wya/3CdpW3/PcUBc6+WK1/XoM1Olo/FyE9SKzHY5txNXKJxw8
yZ8wfAx2mNsxLYLT8VSlIEuNm6O9D66YTZj6efC9QlaeqDJmMmQsCg/5rrg1Io7CuhBvCq8XePnc
lnfHEO9vSCmX0t0vGBCjZAIZ9tv6ICQrTleiGdVBNwfXYARs7ALqz4KfYVZPmuChBNbJig4tK9M1
Efc9tES+rPoJdz5xHx7oBmTW93hmCCtgBpgJUmx+fr37weKui5WIRyuHovtt3oX1P7hUGisgEtk+
6bPcp81zVMa4vRUmjpvVHk+tbN9fhFZpnPIUYU7VbeH+sVPBRg7GbXjBQSbwFYcdlW0nNiN0tSCX
yHFYaNp2W2g4jlgYv0hQHMuhMqWcYGMu4yAl5u44xr0aYxKt9NMObPV+/WJHsBwCVRrbeK1Z7STa
2y03oZLH8pUxh3E6WLSEW/JddsqtE+n1xm9TLb7S2IO1PN/wnaShpIQnjn4BhN/H+5pQx7kuJutU
HBUu+3cxn3i3ldzyucAUaiZkcNgIJJFkxCaXb2huMORMx+hl4qexfJgO7IMqe3PG+aZZVsKGpE/7
Sd5ADm15pbB0fLaAgTnb7jDfpqDBk5O5EriLwf3U1Jt/aNdOynEvxahP5lEX3rc0a8TLnq5lznvM
Ka5EwtZp0j8GQ5fMO50FxOcUlnjjv+4tOqTaFGPx21OO2tctNyNNpQ5xeWMDPnMwFOuUcbwQSyk6
EbExIoWOCQI9CWDtqXXqHFvPdNgkKv9dwmsVJG9HtM4wD5GcH24yUwG/e+N4J7lfD9S8hhvRyJHZ
o375VAKtgVequ94wPidO2JXmnt0s9W46uUS9iEm6r7RXq/YYzjKTU5dRP7+0tYTBNn25r/MGAuey
o3CNhfSQfL8x+rZAftxstDR+si1cLHQqf5iMWubmwT+OR4DZKiKzSPSquaKkBTrXRg0MorTBovCL
5Jgs1fyefMEj2EhDITD4drs3qtOGw+f2kKTqpKsCK+8ZW0NkU0o6wCsh5A/LMxr/mh5dBnYAuYKb
zUSohmq6U37UyMDNZ66Jv2hIIFunvym4jYZBpCqD68UMrlEngNB8dDOFIyB4xdcDBmnLTNZF2lr8
FRxmDz2UA6FmaET6X9QxyY1QRLmrRyg7YqfwrhGkggBYF1BB1nPdWnY5g8o3pg7SU0GZvg4NTGN1
NTVGUjMwpqF3cFuZlmD9otzRij0TwdUC2IgAKu7EBByA9lHGNH/NlZeywyI7KmqLsFj1TO7y8OwB
ExisCwbZY/MgGcMjdm36TFlyuO2jcTUpC+HwpcQ2luwZpMfX1kx4qmum7j/uomI5ZdT8SEcdcc+1
/rS55dGsljQqLajZvG2QD+7+qhA6al1qVeqp6dLUTiz/GWf/1tzOYsaQ8+f5feMWtDqUGKVMdFK4
0r2QjrF/WYDsTECN/Kmmc6Wh86r9b1iQiCVNNDzSMrTDXxqUmZ+HM0gJBR1X2O0zQyPJw0SGRUOj
rylv2lByS0RkagAV2Bw+X1UO2qkWBZ+TsO4kAYLn/wSdBpWfk9e34+bU+XEQueiZ5xU8twdJfA5W
Gkwq4+Dn8s+2R4EV2eNgoWJTAJl3BP/yLILRE4fWxZBteloIAfQuxY6ukPZdZDEb/2HiCUgYxupw
fI6tZTCqDQsVGEPANewLN4t131txiT6dFPw+qt+ZcqOKpsQ4ll2jfn4BWaReGzQZ3n3xwxzF1BzY
NctabIVB2O9iz7NELnnOSPonoVJGIYWZg2pY7Y1WueL8MdT9L/gDgfMq3/ZlOZq6jXSYMcXyXPTP
nzb7G71e7hnmSMZGEr/lxt8xP8Ui7quHqp21rLRqQM+tDj8KFbpqtEae5fB0By6RA0KNOfvI/fIN
+FSGmzv5i7bghm/sVqfhS6ZqO+X+fnO7xhzGKLrCdHfqCoB2P/pRMy79c/HPfAYyOFqvdPkEJAHF
fQB8zphrX4hpgSH2NWlQjJ8rRrh3mrDARabQ+EZ0BhbH2It0dEqKIul88zR17sQ92f4Fm6EI2G8S
Lo+RAgiHkr/4H8tyxKiyXNqU7uUxhWroTjcQtIKWthdKvwFRzTDlVqpAs7aRNFitjOzeDH7SdOKu
2ESCSFkgTj5Lio+Qi32kSP2rOpSQfNyvattbQHkfqXbZs+oK94d9+8uNkiR9pEXRs/Kjh3xdOkAM
DsyD6PkJFIUmO4kc/QOoRJwIgADdq1dM2n2Ajy3nU0tZbJv/tUqNaT9jhLfVzSIqX2o/FTNZRyfQ
G/R790OPsBC51nAya7kZKNCOFtNvj1YgtqedpBVCS2w+yAOlNlYAXJw8ip5M2m6kZ5kkcs+j0nUd
r3qnEhioxg4/4LfKAUvVvcUHuebwgkqOGmpedZAqTqVV5+gXU4ggf540Up9KyznbtXCkRCkb2IlC
j3Bug7QbibY0gcdPn9QDU9ofmYLQRgMmJMOu1PCxnQBHvSlwr8lsCa/08E4AH1MUXJdLy83lYvIR
0t32YA+65uhJknXD1OY4z2dXAhb5l0FlyKHHV3HLIW0+btMxENPiD9hriIiD3SOzfY5/80HllWwa
uv+SaJ37rrXryc7UBXIi2KAmXpkYek7NaKB61KZnLZf37szI12b+SdPnn4sFNu3FpSJko6G2nMN1
1qs99b+ADOPqP6wOY7B2HvQuqcFZcsYkCZBrkObA6oYhNbtEO+6H4uux/0yXooHXusduOzten2em
jkXx3lFqZKJ7gGiSnFAHENE9BW+BGYk4lDViad2tq1H8IHw0dKQSTA5U17dw546GZvCxmcirayLp
l7mFGcoKX3OEmP5PIOmnLfER3jIKoX4+HZvgzy+qi1EvPC9MWYCF5b1aONRAscOFbHfplrmkP2Hc
l479TS044pBQp4wTazakpFOP04GkPTmsxS5ZTypbZLyQt9V1pmehHGOlAZ+U9COwvOlZMMucC58u
6tjDJVNIWofVbQ4QI/4lruMcgdUfgHNmIPtvhT9BiGOdA1Mav55iGtGnuUMcg57IJO9O9QoyeeEw
igBOOnu/kGf0KlBm/3DJ/J+NnZ6ijetYsFbEIOoFD5QK6PFj2oVohsSlosj7vZ7E+5oC9xsWSJF4
iCPn2Vtr2UMsdKWYwsTF+vo78Bq4phI5g/wWnP8/r4cmD+iQ0kfU0qHz2Cusstv9ufDjtmrvAGZy
xDfUk7WswgTkjK8ALfoNAUWepFuUvYphvmYHPqkB1iU3SuF7jnCOTZrDFYrJDoS2D89RAeMAJyQ9
0+tIQsTf+ctriwjeHQFlx7cjnISGzpQ2Y2qElpvD6puKxNN4KIWylUCGXAPXGwHLikkGWpdLPnSq
FgxaHwpdAWm4w3m+hpvjZh52HAR3Vog8G8OwRQnBvFIU6WfVhRglA/wpOhsDPHqbrlritRFN7SKL
pucPq4EVG+ma2+hBhivO+Im3mKd4ei2k/S8n2almCbLsUqjzTO6DC0HotrgMxe5R6Pl6/NCUx+O/
3i4YXwFQHTlP40MUXr+cxhIf39NPAvzgtrqluUhUUN5yTkoQarfF5gPt9kEAh2kGoRDeytHY9E6x
S0ujgziY5EPMPK00o/BMtqjTWN8X4nIaeye5VwRBCwpht+tRXdLerQ1sTG7vPC5GyovaAmL4Uf+r
XQnqjh7bAtthwU9zTXQ88yUOmAFFpFoU/qAydgYpdnsZsHAbF/1ig9pKkSFmuKDac0a9JO7rjOzz
XjLQBqzft6ZfVsrFz3bJBL/l7yHqiDcHqw9N9TNW5oM4bQMcBDYUaUzUOo+UPELpSYtB294iFD5R
ZH8e3lWlANUnyoc31nturPwvyigiSFzAMbhWObAGQ0j/tK+L+dqlejL2+1nBthsweqMuhlKQN3fz
HPTFeaOjYJzs+Z5O9laoGUSphhCqVe5i/ORR3u8x69cobgWlxpWKew7G4VNkbqSLaykCYR7pnPxS
ahV3zeo3ekZNetTLJp+ISzcrg02CwjVq0QXtPr6n9NzXnN4lEOmb7XBtFQk7SPmzT//+6CpUmnLU
+q1sCbIx6sS9ewZfY89gPNeMRyRrRPnFWyJtgtyLyRYPZ/NnmvaClDtTeWHnG3A7zrWo+lLyAPV4
oVL4W8yAd/jF7B872xmor2kJNGHoqNZRs2YNOuH6gvWv+VMvI9xGSlKbDSfHiKXxVOdWmTBT/yuS
qfPUhX7G+qJw41G8d1oWVGKCRGr9sGpKmTPcy+XHLrojJEGZn+SR6PND+jb9YrADuRo9kUSjaQI7
B8V/TihVGcvufiHL0mCYRB/9J6edxVuJx6eWcEq62rL+V9oph1bo5jQcSUOls5j0qkZaLGRHSGJj
zzAzdbkH+tOrC1dxDVeAzR+e8yIHwL3ly5KT2eSm7o0ZSvsLTnfjaVDWCGidbbUWlXx+uxHr92AX
ea6R2x4uureoYJg5Udvf17vlv6Dm7nnkyE9ngboWJo+iQBogkBj4qSUpr0+ssdk4fQGaPE0QNyls
XMbwH+yHHFezgDR71apyhNm6EyovlLixWCVUtF3ngSHy1X6koHXnNA1P4hq3YBsZbFaqOuvAFes1
duMShVNkZns91k4FKQ2gOajh/LIJddVs2YNcrjAujIkKmcOuYAL9fBhcnYcGKMgM0HY5fIVAO9Dm
D9uyr9v9RQIV8fOMRztyNPSTg5ObMA+WeJwKuNtyYi1luSVIFuf7tOr3TaW9NINBIanqjdrSCs0M
L76Ytd43lFbxCgTccxdyPLL0IHSjM5zQXki4Xk5IMHZN5q8HTgU36rIlDcWpSYyhatHk9o0gblXX
0090ReBoRtE4lpK03luNo+O5vEg2tJ1QjFFRQ+QDbvHrwdObW28TrCCg5nlsfPwiIsp2JddbiMBm
1DtZxkgdt39ugch3rBSz6Zg0D9h2mFEvAVjtlV6jzCyNGp2XmCAf5pjfytV+mMj67xoD8icnIVHw
cP0nozBstt80bLqgDnq34OUb8YQgqGC7u4WnhwHL8S41m/hVehUVAEyzC6VgJhSzE8zxga2NPriw
8eTTx9S1WffnAmHk+5uTgH1aUSG+isIvqRpcViQb7Oq/SwJMpA8xpj5Bt4NoEuNnKsoffEGwho/U
FojBJauq2V7JBlDR+Iw3yRaYwId1gH5EfOxnqsHAftflw7iunV5ap+hacH6g3XXe/t2WMMQacBIM
oUvNnKigZOFTGnY0EAezk5rnebYFaSQWw2OWo6wUOEJDHws/CoGvspTXNbx+N6FcDx/CJCgVRaSs
EUIaUwAeBFkToEpYK7mX0DwDObjblUtAD1BebAh+Bki0j4MvHajwgOdhSPWAsNFKh9H68bd+flzv
zMptu+QHVw4K9n9cxqvvLCnwwajVGiMUqqcAi6rkpDcehZGwmUHevMNmdA2iTZcnEbAj7wOLyLX7
eqG9ICEfZgzDvuL4VUr4FapvFor5bsOEAccdw2elbL59rsftBvnaiUSPwAkH3xfFKPZ4+t5EI3Vi
HzgSCjaEyZwH6Zh3QtTGyF1dcqfYRYRgtHUZZwcR5DSvQxp1oW4Wdv59so22x0oa8bJlohZopth4
g66ukCV/vCNDHWKMrpMsRBXoKPPZHD+Qo7AFTamYgOaQvnYO0CQVk6+Xe8glgEwiw2CaFQP/vDnD
GAkIs5zPhP7TT+2q3JXp8VSC+9Oao3QVu4aqVpzA4ZZuRdbo/kGHZC0XOME6LL1UyT+sPlmCMMiW
hTr4gaz1PXdP23CSTYwFnAIwAQ+KxGcxGGOcoPfM/g/IVVq/q03/qPMK8KXQcByV71IIDIw4Vg0H
+LE3IkuaHwr6AyumMcGIU9g5Wbni37qrhfAgjVeQqmVF8w5gOHBzkynenPdUhYdO+noow0kc2TDJ
rIXpg8U1nnRvfbFWkum4LvtvscYpCALgA9f9jL8jhVeBOAq/dgGyu0dDFA+8Fdod6Xvba217wfLm
o8hgstD7mCvF8/JBqtIr21mtuGZvDyswQrbn3yWdHsqUzCq6Sdr9EAqLXm93PDvEXmH+fDrpr2JR
Uu5S4S/Wj4+6bLOsHcR9nxxZ3dE6CyBvGPp02Eeivy0J5ByRaCUKPi5tkf1NXab+hI345g9Dm/lL
IlM+imOoI5Lsbregm5LwuOgzj40Ns0CF9axO+mngL4Y4wYqzSITQl/mtAOwxoN+MvRP6UPtHbojb
dL+B0Ar0svIoVCDWdlF8fcPDXLYZmJWcbr13Iyps7QKt7NCoHIPJ0+9JD6kopoud+OJ5u3TUSJK0
qIxb8aITd8HnKrdFnCptQ4ewL/VdUIW08nXp/KrCSjDmx7x6yHXdqt1QAdPnjbLk++BcsJ0bKOKP
q1lX1g6fnYyRPEvGzY74o8ncjS5JJuz5aXgThaQ7Fxue/FlqRNF/n7bVbbyFjAMI+c74VlY4q1YF
Tv6LN37IbwNiEDTMFtrOK7H8HnYbiRWO2iNroyityWJNY98hHN6oEU9mFv8zQ79GqOFOcjw5Dfmv
JMRoOcx8XkO1GdyaNnvGAGIvSPqA+xu9gOmq3YqoelCXUGQQOoaxpYd23WiaD63udwIZhiYkku87
a1yWEF2aQEfJe18cTDrpBB8bG46139GLQealQL9DR2zonxNzi+CnbX+rttxijr8ygjC9ey6d2t2f
/b6X/yRgNtHC1wcF75KKJewoT9ruTElkULxO+2/waQ/Ik9LKJQL7ZQKlgDqwJ6/NEXmMRxSzy0vu
7G80+r8ZeaMAAcPC1Sh0BSka+OnEPHXBiXiIHtpvUM+oR3HJXKfFcur//GEPDFPwfoLt6+F1Ppc/
JwxJuQCDziBLxAOHmG0f5fPSh231X3cGY887ICjKsz1RARNPWicsEGHYIHOBGwxT+RtpMgX6oPrF
9uj4bbitfSoTqUSDKeAuYTTG4ZthzPgPIzpQ8VgyEjUIMYwbaBffYFF71ReJknZY5xThzNknt3RU
+u7JkHPMX0qoON9pYUBqFgbmYr4l5VcIDLcnycttTHVZ0Gj/nEY95cRVlyPhbkZiU+N22aDaFTYQ
jORLavepElITOnNJYngTshqtKOloEUJXeLvblA0fGmIu9lTa+fS3Iveqs8uR/V0nIN+SUUmwTVUL
riH9lEnlQnMwkhE6H3Gb5ZNviROJ34gFwdIuvRbSo3jAQU8q/P4oP3RgZhhzsT1xrM7q41wQ1zhe
3UV0ZdjkOfhWEmthGXLJRh7ZvSkP4mu53ar3aJYPoqY4e/tSfqk1LlchAd2a/yUCq175velTxfcc
XVM1D77vIxxjh/bZjUkS9t6fqkgu9lv6FstKlcp0WAgbayVXaWNlM9BLTE8X4umBekJ9lyw+fnS2
2QMZrcgx8pqqkeXj6HaKz24cXMUcQ3OMem5A8g87CLE5aRIRpnMUoEGHNWZQ986SqZjiRgR/64R7
c/IRJZTi/9DdSKe+l4o5rLv1snDz07PSO3XcEMYSsCQAX0L9gyI8OYFdvu7hBIeEzd6tFtfoG4pe
/ESuIi7aPMJUb8+Kyt7H/aLEx7Civuod5i3Cezzslddj7fShHZsvutninBQ4Q2XJh23ztLK1Zwaj
8N+1vffnqRbn+Z8yNGYh2u3NAOVAVJEA5gk88qHjwGhWtNEXYZckarsobJrN/FgaNOhHfHfMsW5E
8L22mVeXPpX4LR1xCuA8lyMV7zuFcL1eEirCQ1BgP2q7O+CYYIElUXZDJzlXl2lTMt5EuiFaV3uM
A+EPhnCMKc5NRORqkYvmSdyA6R95jBoGx0IUo4Xn24tYtLOI8x9TOx8JvEKYvF6GQg1PmGTvr2/J
nWtuYLQfx1qhalnbQJnQofT1LhU9j1zFQ54DrIJWtQOL403VIbbGGfZj9YrCHtoKov2jeAUBoqml
4yJWhfD+VmL8+q64OKPUcafkFOl5XVU0osUNW46ctJRukaNUv6EPFWhUVATs3u40uLem9qpXlENm
knWi/nOVnkpM9w3cBmWGtg0H62EIzDTzpokJXk+WXrCJJIWTr7wZCHeT+8i7diCsmOVObWdB/QEc
YD7/AuHsPdQMiTyjz+nzCUsY2uKB8XJCawX5lWo2EoLf/EA2GPDRmZ22RKEZL/ouhIigMI26qNWv
QYBjRABAkH5UGDOb3SEMEN2loV6CwF4+ZKmH4DYofru+tFRtoPvqHG8x4YCABu+uHLoUtHammhWi
r4FiqETdpTA2MIqaEnIHrNft3YPwlh5WwAq6cmz5+qOIHl9EZMypqGSTfnHjw2NhkaHZTJ8MWQoI
9LVOS4EUce4NKK5HvBi7x+bCFl3mxb7DhJur7HXcqNDFFvDrjg3ZPFw14WNAC9cewVHOBOsetJ+A
H+zrLl86KUEP+GD6QKSDuj5rS+Fzof1qx7X5tU0Edg1I/g6klhdF+QjVTCXVWTom0FaLcmkXcHx/
gGQJqoyglGt+7KC78BHojip2Tq6NSZ9zW8DvAYtY2DVNfo0PGheHktePgMnG+6pPlDqpr3vvsXj1
kCVkUB4O1PKDJCCal8qAFL8IxQsEsbip0/RsYDNMSpf3KARnOd8e2xvT8dY68ZJl5SloBZ5BDZDf
d851AqpWYLCxt8ToNyM1kiiHYjhMdShsfViuh5JSUdLaDnpKhLCxlXYhqFp9eYXn7lCvfTqkcszI
TZP+iyHB2Qf6oXazCKzs/2r+QF4EXuyGaEasiu0Yi+Xl89gkCdG/MuIGTai5Wq88J0e9/qpC90Hx
VjvxKsWhkq+kUWWvmFCkuvvkaXz5X4l36paduucQj/piYEX7rEnT4UsoRGGk0FGRyERkNvTs5NW3
shTL+YV4yXaZbF2n3Vcx7icBZqeSbI2zpeGXpR/z4oYC5TiSfJhrbS9M3TdM4Srzq5fUl84uiZTZ
GPnxj4U0yLBA9mpAKYgYhiVu/XdK1wtixxmpyTgE5EhyUDFJwTJ2qiREApPTvTqO92Ra0X6Q4zQQ
/asNXzEdkKbGercX/VovJKeF0ZID8PIrp25I/oRqglW1tp7l6JLlOJhB4mOe3wNgtvvUo0d5t2Ca
XV6TiZKUWSu7HQqprrGaIWI5Dklupw1HAdzrkS+naWOR7rYcW2sKeDEFbPeTdj2t1TAJef8/HOo4
MVcMzBlb2YjsbVFzLuhdR9RTYN75ohoWfn7WPx3WggnikQTliRrvK60S9WcdNlSyv7EqTv0qCCk5
AWpw5L4+onOoYkeGw82QH1gmOSmrkxv9FAkTO07rn2d+TeqspNXFzRO4N+RZX7X6K7ISRwTVhvOj
Nau6EusIcg7s0Lr441YQFTOgpRAGjhWCw5fVI/EUcy7m05HkbsShS+cd4iLPtaxdq76Is+C5OSXl
QnWtMnGVKiErxDsIyhT2olLX8FBzCVbJjJg1oF3rcThBki6uIjDNmJSete9fXgXQP3NrtiWuBWvV
QrquafYQBD4p9vk6nLvFw/5LN1ztqHL2csOQSxcEWnTUgrBbgGCT8Rgf+HS/jUJcPVMNGGW1p10S
L7plec8DtaVi9FhUFJEPNvNTktZoBKux/lhBIx7EQY3LgnZHyAzeHHi0A7sao1R0Q2fkOwXnOdTR
ER0iIGvnodVUwNYut0eTsidGHqb1CccXdMdCxZWxDF5d5G/MytfGmpaQHeFBHYe5ufo4mvxqGIB6
xBReyUTQdLE/vaT4UsE9Lg8qV1/2cf1btsHyVw/lTOooMQuCfIYOE57r5P4H7CxSmrYniNtOJmzA
eRT48iEgw0ilnKHpxQCpvlt7HeVWKKA9NSglcKn8fRHOOh+u6PKUbVAcV59BV0j+2mqiN4NydRSj
RcHhcMaMmXgg43tJAi1+itKcyhynMuEzOKTwj0ICOk+mI1CD10GSrL0pioG10JpZ0HhhfVpgYeVG
Kq5cUOmFJFn0juyA+FFGiuPLBbdD+isgmce2pDvu/BWrhlKxM23C3Un7JB8ET2Lorov2DqCP8zWQ
KSg0qUXoxI9L8upuFmXodk6KzrDbq/15mR7YohSGVHA0/rWKbZggsgftaHcfI+F5jAcALVPAyjGz
8pztfX1vLfs2uPZrJoM+xdEbcEATSIDxbitfImeePLujv2rBbMCDV2LR0qfUrz0OJhuTjgAq8qPx
niawAvhmDzqFFq6rlnrMtJ2qVognCSHKYlDGXo6lpnEPxUjxuuUgpJG5chvfK3WGHFu5IsdhOzlc
DY6dgeWKevCxzklgPqX7BiWatyPDi3CcWJFv0z5+Lvt0TW4w4HmrpkXSqlTomlpGei90szAlkG/I
mib7EfB2vq+TmZkMYlLgaP6XOUfiiTIaLn/R5Z71VmitMNHyii//w4hcSEaNg6K7WeeyLwEPImLB
TE9Dl+J0SUAX/0didl1voQxN2zghGClH8tVyZiQeTBe2Y9OtNiKwz7xP+7Bd4tVUpreeIe8Wrg+u
fUqlIiATW1sphA1prRKrFHgR6cAc6CYqNs3h2vI9KJFs8m5gQOf8y4c2u2VmJ2T587Rk3ShCWysS
CfGlhkELmo0XSgvzmVpNN8o3mgqA1iefMkfS4fgpA+xRt0DDu4OXdtbGXskUWK3TUFHqKHX5XGgD
Gnchu35soWYb4HnT00nZjyu1MJdDtWbUKG2cl3efSJsrW+KqA2ONxQ+OJy7WM9o0IOJ9jgbFbcz6
pwn5aagWFdTJJCCiV2E9wLjCp35tZSTgKWXVK8U0gFLrPvUbDBnC/VE37CcOapxlDB1eK1fQN4KP
aW0LQZiaQXuvye+ERTeGjAkAYFMU796fT4u909EcAoxM572Ay8TGPpo2xMXmFTaOCLnGZLtOogZZ
7cd1fDAXdv5LzcxloJuaVxwc37pWteHOsHQBoWq+QozAy+IuEIUK0Nk3+H5VZy84Lx9hmib7k8Qc
Yc4r+ap7mwoOToet/L1+fGM2uxe56DUEwHU6lyeZ7WWdtHB7ZEZpY5kXyrUwewOrGa/PDZRuYn4G
rQhjrC6RDJxj1/Pj1Q4XNIlWFfibFhem6iXETYET9Cfd+V11NOHQ2xaS/4iu+4XUBmWZMKHF56Ul
32TbTI+WzBxeb7ocYr/CzGJmBMANDttRULxW72vbWdKq2nqcj7XGXo9IO4RGrYk5rT2rNwK1bqX1
3bIB/61Xz7H8RIrcuKXuSRxVYjEF7bGvWsGSga+ZTThEbghDwwZgakQItol/9eaS58CQxsw/bGoH
WwdzojJq5jDtU7jLyiDH1Le9zK3StW3RT3Wpd0nZ7BfkzmLsB+dticUCNvE7X6J6OXcoRc8FWScj
ImxtRHwQR2wm5k6YcYX/WV4+O0fLyjlb9BQcckwFAJgubzw0+LgqwSxmNHD0/Xp412SQZeRtvwpH
6aYtO24SPzj6pDHy8f2d6Xd4FSCp5SubVScicLToeKTmj5b6eoHMtYT7WGYr/dpUZce5+igcz+xV
/nPkjxnX9T0uIvcQc9q9gvTbKXuMvodV5wdXNM0zAqosFCjqLGGR12KGRjJ8btsgYvtxeOV/k0WR
lE19Rlja4j2JpECwLk1+Z5ArA4fP1hvK2sQSaxZSwOzWA6KbNpmesJ+Ob6elO6r6mDLXM3+UBJGw
T56uLWvxLsV1GsjeW2kiChjUcW5ydKbvm9MVxRRVmoyh+HcEdPOizuh7/KPBLkII63KhHyx8bcD5
qH7CK41DRi2YUPsERcurQE2CPqKtPpFln6ZPsuCzkfmwXu064amarXk5PMTuFcCzGcTAfD/yT59t
sLjVvsycOd1p0Z5cuZpz+NQNzwwTVl6yCxueGWA7XQUaAiZSSrGNU+6G7IninqAq2VXtteW1tjj5
WyZaSfFLGRlLmVON9ux16d0wqUUM0oHFnfY6AmtjE5Q0VqCtODvdoors2NuHLrIkwkfSKlhYe61q
/6tK3C0FU3yHa9aqJCV635/HxIVTvdXWHiffNtk15xj+d40BhLx0cd3omI6gbPqgqfa+7t9GsA0W
8OY2yoPXdvXglFgFfa2Yyr6RFScOP4G1P2GYO56RMrLHoCJJ6qNqMBUNH3rqULF0e6O6l22J891S
Inr94FfsGYhQLcwJPIg4kIWudVv+ydx6AWRCH/tzzIbZV1XZg/913R/5X2tkgVRqaPQceSSHSF2a
Pb3wQOx8i5K8WJmtT6gHL1rrLjTjCtRmorQIDoTFBGo9oi84LOQmIKF6ArObB+t+Fht1L1z+T6Zp
bHSnAxJ41JUfrlJbJ381tvz5G6IzHFxDKgSSdsgfoH1wnQAV+Y9aL9piztLPqkVlIjGnTHjfxl/b
nJZGGLbqQf0nb2cBbScILf+5Gnhpbn3VC6BY/Y6IrFrDiwl9RH7wzXhgBfJVcqjvFqMkqZlGZIhM
966tt948G3ALlYCGMrPK3KN1WnHayP5F13t3FMf6VyvP9z0e3Tr0ccHdZvlSRooLGlOHotkc5HpC
Z982N58zM2lgg1aLKFEYvdbUAbI7pe4f9UjRkD00phx0kvr3vDZaRMeYij2kF/LCRlXwuap8Ip/K
pQAcRFhZMh3sS0FcftCCrbBpRVWhyuExS1KrzJ1yy7u5be5hzGnFOqCHNYcEUxJFrgFaXJrMdPHf
EtUmJGQ6OKKPWDjFIJD1c/Deq86rQH2/etqGJhiHMNv7RWXLX82w6GpymcKq/vOX/QVh/EouujD5
Q86YDA30UdAyzPPENzs+wP1d4MKnE1++Y7QQaurjGabAR0r0ZAwhzy/IcTSZbQemxGaf3oTJtjJr
ss+qSviILrErM8AmWaScggoJQU910PESEzTkFSnWhlc/8EDqvF5WZqIjnit5GfX7iy1YUj1edVNd
1fpiCPXJnmjQrOsHyqfa9Mh5rGMVt7Mp/6QzG+LhZydOKstVWH7fswnzmZ2Y1Tm33SUkcag6iE66
ufJiQGaM0ZMBpCfMBIR3tgo0TNoxVwz4Fgaooeb32riNsNoziYDYuRYCjN2h5HYNjXuZbRbwlpGI
pxyvEZbYra66cILMH7f4OeOWJEZUPn0iU9Qik68VSGnQQ62VJ2VaB5I5+H8d3RIwzR5XmhrKOKpo
TL6bFTwrIQPpRF88ApMhRUShbWPENMhypoBIpaCIPGx1dYG8jOnNfEx4JWaacQAItQMdYd+eHguq
T2bWqfjwJIoNykIVzpgj/QHe/3571yp54J/578WGCZNVgrVLmqPQydmesxhgwIFrEyJKahhV1ru5
XC3+G8umTo3KKsd3Tsc5tPL2Ax+i5yyYPtMav4DqhkTRhqjpJ1fT28J+y7AJ5a2FTavimJvtbKEP
V97vu8y0FQUfmzCpKMR5cObvHIa7tHyaLHiD+fBAP71ffpT6BpHX3mzh7LjywdBMNT5FXdVcle1N
VQ2nP9/yKtRf4gVAgpIcTiGvb36v2vXdD95BrjUDr82nUSrKrgJksYQ4FEguTZDl6+TDjsilqUCl
1eMEEGNjY3AmE5lm3XRyjcwb6AdT2xh5u6k8jxK8gqbuGHP7ZzCIYLaskN3yQVJXkceqnx5ADHAV
lOglrPPwZhlBknxMZu+e9tPDQGa8GXestZCi+mzMRoz6HtygeI5K8CY1k14fzoKyWIIV1noQS3kn
/0oihBQ69jCdqGbzzu3zPvlwbficC+82VMOpwPkFGdJ7/tBD7GhkwxZcu1Nf1sbRfEvsm6VnKVvP
ivqc3eRbxPB3opEajD92xTpPOEI0Aiiz50z4au4DEmfTVcuUTrZqcmgMY76yCz/vCc1Kr+vHZymo
ooJR7c4z9swxOg8LAAYMMKf6JY3Vi1j/mfbSdYh122RXIofXgo10Hs2dVMfB+mBJ8Ae1f5w8dEVD
wxE0E2W/ANKJ/hw00U781GiAPD3GrxZO2/ZDT/Ni1D/qk9bC0S7MjZUVVIn6jPhd7UGNXK1tO1BT
vkvrMVaQWajFzshCXDRtAYCepXMuMF3HPrAdUyKi06jIHbpiyxwoW/swqNNnveo/FPBGFIGAOitM
ZhRHTcU3WyNggh9+NSF2ACNhuoOCM1OqU2k1qS+k0RVniXxSKQLH+vhgdJIZrojUCzbKzggsWEyQ
5pIQcXJYsuugnJlthA+ZNhfJqB8432IM+z+FPUqlsS4///VvWcO/vjLiUfFZbZK/bLy+/Uepxygq
s5TDM+Geqz82yECDVAYgRQJ2dGLGQi1Ywu9P0CN3svcNmOxD1CthdGnChDorP+GKXM8l+KbIcvKJ
umjhmGO+BOwnzXVYy1aKlZwK6USKHdA2DLZGPjSt5dxQ3geyFQj+6/TnwEllV2jmXBhRe3gRqJK7
ZdJAyxCXo65v+TiK2GiO0B5D26Peq1eccbu9o6L5P8UDS2EGFl0202U9jC6/+NtcaBTXk4U/8THw
7efUKQhVEG6m0fCBWE5mOhp+WSK4JlJWhLX7tWFWBn+LONaFZ8wUFA9geVc4XcWWFgdvJ1oMlQun
XD0PBxERdA5n9yTrNY624JLLaGa+iSYMXrKn/qBb8mbc/FjIQjjwkj6ytGCIKpyIXMFrKtLXOWKU
7YeAHkCGryQVLaVFMi3loa2lcDPJB/xanCr9O8JnnuJM/O4j4g6/2AGslzjNXmvFlOIw24wtTK3i
rVwcFRfXNXtCCA4nzjxKjnRRUMxY42H8nQL0N7ogRrRWUCnyHhb1yzN1SlpV8+T+ekpkkTxtfdSY
IoHeVZsNK6C9rdlfFUm13ZaOMJ1TyxzF1TwTb7HPpRtyA59hTBaxKkPiYyrL3Q06/CsS3AG6aQc+
wX9v+2faAT4+Q9FTmvfYoIn+NLTDPo7G2cvFqnRByDlNla5iGubONItKn60H4Ums2kSdC7UXI/xT
+pI4Tn+wlfY7JRjbD7o005P7L7uD5UXadJrnywEvu/zR/cFPFT/OW3lFpDs4zpzyM5LpXu5UUT7N
EYFc70FmG64H5WcjMcXdVtsLc0z2EuHLJXS0S6KdBL/Y3SHLKjblI2jwkgl+fsmBeme25djNfqR8
tCEKGBq9WLoNPixuSAhBXls4sLqR3/yiJsYwsOD/JF/rMA+cHGw196vEMMtpICCRwek1nrU9CRab
ZDrHjXnCrS0vXnvddR/b+bFTobJzxVklgWHtlLfVwIE0hJyvIwSi8XfNwiu4lDtQX7Xl4dfdIITZ
3ETVsy+9hLYnegYlEqu0wnmG4A9UjIbq2xP3lzot4nVi1vjTOAb0FrQDq7nQtgDJfDy5dHJuZR1F
qF9QZiwKg5TtZOfQ/NS+Ryzl48XJUeBcgZk3FQcvn8c+LFJZtdMX2Nwm8f9rYbpNaGLqT4xla7jj
p8UB93GunnwM+yovma+4Tua1AmOux2yq79LVqC0K3PS7UkOq9OA03Qrdxbdgq/7tqM3IjfEBeRrl
mNgk/DJ3J4eSk/UTJYkOTXHJK+gmAUc1m/gGBfurLKzvhaA1r/Ns0lOxVAtlfVTv7gP9CxjxbVro
qtOe49CqzCN/rQbTMAVmsQNh1QJuw4Bggch627gVQD0DAitVUV6gs0iNM+/OLFLbG+NA9T7Pe8A+
l6qeBKuf2+m0JM5aqO47G9p8pOdT3AydoSsm6dhkLmGjOb/VeSIN4p5qyW+vTtcMLJIg/tdri6F2
Z3m6MjPJcDt5phT0vX0IfJHiqMmiUrdh/jAN63ZalSX4/UDTLhQ7YP/k1RCdahEGgWNkxhxUAIry
1Mx2D2heCPFXNQqepkot+HXEP4nqGzB2V3MQeKFM7CG/1JsIEifJ3WDuatmciKhEkL9DXTb20DM2
3qU7YKBHKbmWVzh5b6QlvRptF1Rm5WAUjnl04lKK9TzB23aZ+rTVmCLAdGUCI0c0EKLTN9Qf5Rn1
J85ECK3jyWyPyA3/WzAOSaoDDDq5eJgGba/pg6X8UJCcdxS7OhmrSroLfva5Oi2mSM+B3m0NTxEr
OlKDzlp5rtgQjoIwe3JcpdBfyxI8MT2Q+xP5+oQBmXy1XOGyplDa5Nqw11jCGEKQs6PAXZd60KGE
e3AaCExtRVg+2dKVkbVnbfrXTbm+KVdFcJyD/D+KIEvzybN5WFSaUEnAsa9bzfSjmQOC+vIDB8al
SX3Ewpypt/n14uzMBi5g+F4+3kBSYsbAb7wjaspLyuXa5NqDtCt6V2WWfBqMONXzTwSjvAenxEZN
ubVryyT8Ck5miVNSj9PoVHxU1akue0mAX3HheAY1doPDPn3ztu4OEJIWdLvdkIGR0stTi4aLp+jH
9YadiMXtfxsW7663UuzlCOdj2SWnrdHIwsuY0sVGniXH/vtBTU43i+wow6Z7tYp3/PZozx5PjBOx
KuMtr5+JJXGyXncuzAnwfV1ncGkT7hswj8KvK+mBkMIVIUSTs3gKy7hkMxIDv8OoRkcrOCsje+eg
eIptdDpetxHJ9nZg4N0rF4Ziit5gK0e/LEemq0/FUnkc7xyvsIrElHQn1BYyRewNDG3W5JDfq8vI
GOIJ0bwR5q8DlRvOXbqZ1s3MilrQ8h6Ot+DK5/S9kACQz2ipVKVE2BrFI0YCyC5wuiqUuEu5mpjv
D/fVq3cRY8bMgRlYq+PZ4+tQYCz6zdi877P6DlqLvy6iW/6XDXuiWj+x7STdANlDkTiGptXsOKu6
JtiC2A2kxj/SDnOkc/lf5vWrQTbcdd92PdbbbJFBSY7XwNU+slSEQbGooXtiuF5UF341BofHSMBc
qMGJzyzQs1Fi10ylbSxJGboBuaZbXSKIhLmdGodIeblbrqdsu3GNYK3548QWje6Qwl4otdnPmAVK
6iEBAFlb4QyesuUV9P94bCnQJIeLpD8iOBe0c2c3vl+Rvg3uuBZ1xzdbnxGVaB85LZKtU2CaBKBa
xeAFcnHobp6PfquT01N0qeywng2cLFAQxhlURfAuqtbq0LAQgsgQ8te22+erTnXjvN9giGrv9gjT
USHT/i7LX40xoGZYUrzpk4PAfEe3TcpGmcdycFEOllTWi0esj6xoe65wNl+gWVZTSj83K25eTtff
XVxNFQlhyaEahiW4/o738XkRhsiDklGg3IifmMzk2Ip7mpn17sm0tB18JyaVOyK3If9Miq10nPE5
NvCjWo9mx5CefqQpfrOd/oDeqQuZmE6Aj7VbA4m5U9E02BH4A1H6tEK5ovp3YER98weCkXmYwpYj
XensOt1XsRYj/8w10Z0clvZterp3BZ2k14d9Ss3MPb77QgzlamlCsb4stsd84EiTSXRewn1PHRWw
dozOeOx+iomVgn3DuSv+hhNvzERxXSZZib+6Jl6NSKL54qmQtPc1Clb3Bix+HjLcIzyAQyrtYN2g
IjO9uPZBiqe7ckGVrFPmKiZ8n8idYZ198W2I4Fg3HxFYyyXyJFt+sD9YigE6mk18yPTfh3t9Xvjd
jX0+8G95BI0Nhiwe4GzVohN+Nh19QcDVo3ytsbIyqed5sO29IwzpF7LL+vj8zBeMJuo3+Q1qF/d9
gwogHHVlj5B08HuO3zVN+9Gr8YTp/nj5Dgls+9k81tGLvFeKWEgIGuUzIGYCpWqYlHOlvEj5Swaj
VBwfN2jteDTQKL4ZRFHBI0j4sTNY7B0rEYxRLZGSpaIsbFDmpGPrKy4n6F8/j2HsMWYu6DaxwekH
JHpYj0eFs3nZY94CNlFeV/LcbLZSIR/rKk+w8lftLmBEqeHyN2xHz6O+FWLlHV/oPV0lGVzWREzL
zK0ucvoDxStFvRrwV2B55hh4THAU5KYAidVgOmlzOlhMZgvA8F02x0pgk1YtIL6AbmpKW0CCjn2Y
q8AKewD2BESKIRTwepaCNxnrFa275k9dclV1z6UiClXYpOtANQ8c7tYKwHZyh3ixroOeGYh2GiGF
5wzWEZjAvIzYi61yDimRcbOj2ff+F3E7ZDCjo8OK23ge/GaXum7KFGuh2moPmFR2Z/C5RpHstOk8
TwKlij1yR0MxKbL+tu5E5zOfmvD16TjFDwvsR69VYnfCfbLkQuCIY3oP1AnZ2vaxh1N0g6bnaZny
J6nodnbnz7pT8DN/raT26BRZhWI0c+GwctcMNyfQNLy/1hyyRHou2TYiLox4ld+B7p2pJ5AOuVoA
s2PqG4Sq+D4MvfXDKAAUOFx4rS0R7OEfi4Z1haPMNlOPk9BXLrVuxF9KeJ4CH6zXIUozlPpKZ/Tc
f3ZPX1heX1J70VuB5FZ2xPWOIjYEhy6T2gKohTng5KPya9HYz/YfwONG9fBfs3fTPCy5v0hVKmsV
W1Ia7vmiBjSkxoGLclnzVaeUTlXxYMD3e799BJi/Cel/Y5t5WTUpTW/6Y1SM63kgFTD27fFWmG6x
YJniXwGjgV3lsTdziabHfb5CUkWFYK2Tomni/oDD9RnjqP0XeQ0u/HDqu/vxULDVpttvnu8OFO/8
ptRAB2pcny6JTgKwulPgf0tzPP07Wz/6sPk0T6qLqqQ7Xv71EZEsxQyHibjNicVvfs5SJYXY7fiA
WqLloVQUQ55JViPkA/WXQUEzKT7Axc29eaLVfZ8E2yCVCly5iUYy6kbzhGoEp0vVsj4e3QoA6s/t
yEJMDbrHts88J4wYBEyGhX7SSuEq2x7/Lg+LbmOwGMsSTWg4xgvzf2X/halH1Kzx24lYtJyeE9mt
mBLFEdbV4CIPA9ssRz9PVL79Hx72n/5UQ3pnrbKGpE08d0FUZp/M1Wil9wjf2cQknHs8CJtuO3sd
pB13QW+68gWvipX1Yz+a2zZZcxiCMguYQ40ns37KJ+f2HgxyKydRCPe2PWKNQReUlvfy2Nf743Eu
DPwtJ7f2/ht3K7+tiAc5grf5qO2/N96TQhd7jXOVvCyyrMwyHSPGvEiF2edxL2k1LASCbTntFaNW
OG7eCWx2OjpbkRmSrk+kQCJySpXyUvaZ4Lx1mHGtZlgH96PsvWUGZGD1xuD2Ye9YmTmop+Ws1nOR
V8kFTwJRnDai5V/Ixm6xx0e0SMlEk8K7w6eGEhQInvSBFcCRw4PVCF7sdMVc6EZ25vmwNWv4Q4QJ
IfDC87aRqUnFNT8Lco3jo1XBymzviczqkaq4/X70VXzll6ICZ3drdhoWluGPEI++auMN2XPWwNJi
Zs1dPfqOo7cT0mFgb1SoqdiN2HDKeWI46heGj1ZIx4U/BMOVi4Cr4IQ/yt7Wgoh5wWaJyShSV+19
/GZc7vORKl2f9GKPzc0UFVPMUdzxRioJ/oo4FgFSXWZy3OFpYuz8BJlDAE8IpKzPAFHSg1UcPjdU
wCes+bppRhSOjIqK5NBy1RtivyzthJ+POORedFt2JqJGKyOngLBKzSBsWMdCRKuMPhOyOJBASmOM
IpqA+9eMWKhD2AgfyGy4+zwZIlIfCnVlVZka9x6+RuOZtXsicBenWHKllCPnrH1kWY/0hV+wBERU
SNJ9ZcwQfcTPAabclsjE9byR3x5MYCbbdZUOKXDSe/dtywWFoYhSTDlesRmuhGBE5/JiOJzkvCEN
9DZ2jw9tmRk57YlHATkqStvDKN69dA0oppDGUvf/eH8UsfRLduWV56KVIepQKgtiPhr0C9AJ9wbI
Yr9ztmINkgo2tb4PMtPWvLt2yUr2ICKSFjK0bfrHsFKbOFkzNilbGTOkVoubyGT5EjQnnIBzrmXA
LvzxNDvazwmgHv9PhbgYJJUskEcEQJgV/uk+Jw94b3HyLZX1eOE3xLNmgyoRkkfjN+Ym+dLQ0Ov7
PLxs/0oAa6YxXlHb242Nq1BzcXHv+o51dgwVasUmpk2f9ugZBS6TcrNKh2NCtXrW+eizNLftIQRh
kajS7oJw+5s4ryTDCXYZmk460HMiAt9fzp9RcoWRToY18Sps+7+9z1W51obeYb3vsOgzxvskMC+i
Z8KoY1LvaRPfOc5WM3q5wydePcCPQy5zSO3q7bq65QpM04g/8aWqNSLXKsqlF6A4dU914F/u/eRG
Clv5P56PEum5eEtjHXcoZDsVg+q5ltFbyv+BqxJNRdhcRCgLjaEi9gbaEFxygalJeY/9p+jCVGib
+q3qgUzFc9JzRLWzSo7ZQqFi8GH8/Tu9Eo2yuYmt+TDkgJn/2nlG7YTznT1nY04S7DuBvO9bSZwn
zEr+Zof+RzEJRdGoM4gasujEknNamrAE5bvbNpHrwx0/LEeTTjelbtfc+Zi7VQojFYkrDZMtXt5E
VUkgYe/vzeeMFRlQqB5tu/zZP5fAJ9bzrKsLtyNvuQvUeCzP+tzQLfXwlPRmlOZiab6aFYF0KNfB
DJySdHGEm1Q/kV9Jw8o3njg12hrQYAwKx9TLW7jaCNlWgJ+ysAta5zNvUNBFD3q/5EDZIqa3D5sP
3KNWRc0PCEWNMzOxAnmIXhztTb7VygjcRo6q8bpbDT0bh6mYLdkD6G+w12RYi4Dx4491ruUdMOh/
f8ox9et4dHzGfeC5lGBX0QU8V2TZmv54dnA7ELwVSUMpRMikq8e8mAdQ1fbNfGwWhFG9jGw/qYwv
hxc7cK5+p3EbpA6YD/W2KYIoC/b1EtuvpUImypTavLEGex4khk/gpUGeiQINJY6Gcyh3jKaHzagE
n4LBPbqO2MV50DuFjnOl1+BHe4vQZJ4fEBD6CiU55u3q0HnEacRoyqf9ZY6AYFV/yI+M4pDQtQak
JGkCVH7T9YkCJjyF/KH4YJHIOMpUhoDUpWrqrH6AYrEWVZhpE2MvrVk6I56jPbKDZ7IRmwQ5/Gld
3Z0PcXpGh7koGlplII1gahzLcqTlA3n+Ixkzc4MVWo2dWro+Eo6MebigDuYrD5CIMOrnWs0iwvmF
MnUrYDbOGwLDt7IBhRS1YRUey7PKZLKzW0Acnm5bH2P/13JzGq/w+toebubDCGog1ZL+UmEhh32I
LK7b3ap860WjJ+PAFas46ut296ODmkmKkvesrqHM3BQxgug1VbrvHump61eAPQMiwwTNR8LI7wJJ
th5kKve6j0NRLV6u5i803fT+RPBtbonlk08XZCv42NjDuEzmMR53pMUrGSN8IA1QxFJPDEUYCOgE
9nWWuF/4grSczyofyetYf6PAQVx8lNly6J1vBA6uKSaSL993WW7isKaSafa2qWFiGQjLSk0SwMov
jaLFL4gLQq8Yr1WWVeq3Y48x5iDMhWgIs5rizz6ZdxHq9O/oRnvOklCfK8xwl8K4P0C3tQS3m1uk
jrTyMk8InKNxUe20D6xEe9LVXcKhHBpsg7FUkk4P4aIuTbt62qtfek3f8tTdn7+mpSlvGkXuB64b
wpD1t0lTX7+Q0zCMl3Nak6cypvC4mtQOX/vb7eBZ3KQ9I/3USorUMG9Y5t5YKTE2mGtU8JOcGswt
2qWZXXQz/Bj6fTZnh5rMXWdQhDwJA1SLVBmtLp4bxX8oY/JchgivfwHZf+HnOoYqWSTCgp0Bs9KW
LRXb2sthBhC8nEgpsFnVPBKMTNFJHFT/tI6ZbqX6BSXs3csKUNkE4QALPeGioFlpx6/hCP2CnTCZ
SAzLsKzrBeUyiyKckYJHt5xqahb0RzUcR5XoCKp6vhONXNjUUEnUsRn8+zvX5LG2ZupxZiDEvSWu
v3IoNPGT1FFTHZt7A9AfxF4Cf6xePuMwNXIuHeHyTImibmUWFmvzKyFKq6gB42oW2XKgPvmRXqxK
ZnNN56geiYxh2g13n+CJ3LjJ0pN1F30uZewLIcj/UPz4hdlNq+JgrHkJ+8xINUS/bsnwSpH0GP41
68HC5lOtDFNBTYHqXvf3S+MugeFSYGAC0yncq/Wut02Mosy9VjLp6NbLV4KdG6u4xRvLwvT85G4l
EfynqylE9R46vs8BisZRaL1mPuxvhXU7QnYmd+8dq1A+pF6Md2i2Kq6hg80sAYMOnwtQF1WvEPMk
551toBBqOITtWeKWN2t2yWAzaGBNXIGlwA1ZlVYe11U0/pckkGNg4bBdsS55PEX4Pjkzp3Nhqd2/
i3S2d6sBf+zgSTAJnA8RzWXRx5fU6Hl7c1r6EatUvdrFLkeLnwnQgNs4yUJUg2mWlItznc6yU+9Y
eOGn1zesnd4CYLLO6Tweu3jgtoU680sU9NhmfAcuZv0mK6mexoDoo01D9se1GgzMOdXK+Ffz4FRq
VMalZsvfGN28cQaU6cuRHcaZ9BrB5ABcMHIH2StUz1R3nu6Ju4gtmNDRjLoAOaBMdFc3acGHhcRd
JVO5NtDDW2oFXrAQGPqLG2aMWgQI2z5L+48+x3m1vt/N8jEHvLcAKkCzPCstS5bGOZ8ESU9jeBvD
LLj+KG+DpRHfTHpimvd2m34B0qG48qGIT+sw8l5ak3Qf/SqWhQBtrMtmtwbH60fRUe/4imui3u3L
O3c88QoBbuNMnfL03ahb9o9/qbXJ7bv6Lr4KLHhnap6tItC3SWr4X7adaTlsET/Dxfd+knqolbsl
tNpnEWHf97Y/mldD1F3ke+8cg3g2UXqORRV4XL1QhTe4gugzUumPZ/HLxWh6Bcz7BIBwCdu8lopM
BPZEKq1tqDHvIsPif+QzjobEJcJet0d79YncKE8paj4ceBEQ55lRyPKVfATzZ5zmKiipg6guiZAb
38cw/xH9Khu9BxmqPNSA8HKd/gbva4pFnQfyVnTGx+25TvatppZggocaf2UwrZtjKWvw7mtO1Rzz
mKNwXfOSlcmt1nYRHYpxRtN3762te1a6cy9WlmoM7+mtlieLbP3FMsRV1PdXQt3OV8aVjKPR3NAV
fidoUNAoKfCZ45TD1QGPgaWStvjujKKems8ykKhawqEV2NIcaVq8J/E8WVu3S1WxAfgY5tm8Unuv
yPtC0NE+UdI/5pE0AIN7R4Q9gxokwy4ZXZ3R3Te70VoiXsjoQlD4aQROg91KmB64s07pCQDggCQM
uQKlW8gU80+SOhsVlZV4ebYuiCbAZBhC822IQYAfZ4Ck/ZGb6IL9FPWTXST21hJX5uy/Mi/U7QlC
KEmy+vbzh/Ppshjl/qcE7azsSOphf4F9b0Licxz1j28Lwpwg6dzElkBHymewKNQAqt7wbFETR5YA
jpmt5hjgEkboUmnKQkBVCSGh/tqFmMTIMIhof/AkZO531BtdQI0Jx3IDGB+K5dbJKgPuG0iFhhQq
7pWGozNMUh3BscAxbWcA5GEDi6yJi4279lPgs1NvCvZBFFGOcOccA7cy73Z7wt+Cd05mLqi2x6xV
4fWx2CoB0wf0jUGVPTsFI84gXjibyovpzdT9hhAQAJbrZ9/bui89TUVl5VsqDDRMNQnEeU0p8Bwz
zuq/n7e4f9ZT7rmIJE6OMfMOxzAEFTs51Gkl7rDfE/pFl7O2XUYWjuGhzp8K3CQ00v5tF+Z2H4oR
RYkZUrCCqjEuC50rPoIrRG52bsYACVEPk/2rvmgpf/BSthzzzXO0p7VXvCMTs01mrwQaJMLsJhOV
luELXhg69cmCMi1wxtARu0wbrLXG2Ekp+fEv3jD15p2z9jNvfPkYZItA68+l0MIrHFZYdHTJbF+d
GHPSsFWuQ9ox3kerM47YkcWKkk9mpu5zxSjGuni+59cVjoZHBMvoW1vTxz+xJ/Bv173j8kx7t7Lz
qbeI9q4K5jVUqFa4cK/Y5Ea56jPoJwUXwgKs1VhcGX+h89Wqa60oyV0BWiwc/Ab+FYoHKrlh3jDo
mU385rW1V6GKQitjVz4PV/J1mYwlkSdkhTIWOPi1716fLu0pXfpNzUKbLfsC8ScKZhJDa4+3SW4g
3Yhz9VngONvbJJR28qW9qTHI1MoqEfwOZzdFaLQ7i6V+r6HaA+LDTMJXwZTfGPsFl46ASKW4arVt
cBQbsJeVDMetGOZs9bwNykJsgDnnRr+52S9WAdNHhcspivqpR0Bv8TbRqmJVNXFFJZ4J7nL5I4fL
jUrZmAgmnVdVSIYyJIEK1Kbm/n3RQBhoJRITKPrHX7Ljc1qneT3qQeqIvzxhx2SpID4g/G/UtP+l
puSC3cc991+M2l/JpDMQDm3t6jMGYiex8eFe4eFUZCV8TrokEs8qtRcfuaN1d02sGj6qgLdBbw+V
jWUglkUM2SIRYHb8tfLCzNw0qyeDCaPqcaxcDnAZrPdjNG4xBdCcQHYY7PVXm+wdGw3OX5rxw1F7
k2q99WFIc29hk50IqHONk32iBopTEG3EnYH6QW3sec2ucRMdPhRr8/45Lq4YtiZpZO5+8IMnb/XX
ikLZwpogqa+7JmSWx2mBbOO53xZBS2u82wciy9Z87lq0t1/YYoO69/dS3jY4hVDHpq0LZdat1HWf
QT9lzUA2JolWizC8juBEare/A2asXa3yFmnb7MhjYPlXmJMDBJQZ56koT9ohhYar77W8irmcb3T8
Ez8zl0EgeSbgnkYKOg18pxwuKoF26NkhrmF+ucWUl8WUf44d4qbRy4uyKPVmq0Msk/e9pUX87suh
/Bul5K9eSMoGRsFf74/FN/4r4oZJL1WmJjBs7Wn07/5sqrGdoPGhynjeohdR0j8SBN4vjiIucX8Q
gEOrsIZv7uOI8voxLEy5DIPC/h2I5XCYuiq20CnILjWY5JWIiWym1YRxdxjpcDWTWcahD5Iae2SW
mSLcGFM5+2/Nbqb6sAzD5eJ/hyBvzb5Ov/KcCfzp1SgBZ275mRf4yotAdIepMnh5VRBb9TMmsMFC
XZMKi4T/p6SdGFhLNYBPAV7Cro69YaruuuJGdoYRjK2ZxTMiNVLKF1Uk86tPxdVR2xp5cvR9GfjX
2lTobrj/CtelDCGm34F/ApoSv9guXXTvZeiLEm612ofaZpumfDC0LsaR7xkw+pk+HPChhHjiG8DN
ryg+qgu6AzBokcEKAhLKca29x1rSdIFeZWicZUIJfLuERcPX9ymfVawFKylQ5HixJZ+t/tI3HGWN
xs4OzmFzpqqxOPYwq4R0mcGCkxUTJ81HMoUi8NKv408ja6bI2qu9KWFzkFJkVhDBn2mRxynMBPw9
+KtxsOPQeZggM2Pu/v5wAFiM3/fyrdEUXRXFaGcAxHITxALb6LAZkDEHzwmFQXJvM7ni/LNmpKJa
Jav+GNCMDz0OcoCpyUMuuBiSNwOdbDW2CaOk/fhsTWZei7lpggc/e/GdHyVfAwOHvy+EqshckBOq
GFP4JNKC6fwbyBtrKJlk35xzJl365hk+SN4PPrOb75QHEie5VvLvz2mKHzeXn8m6EBMGy8xn1CZE
/R4F1qZBOIIiFd7sOKbZ+ZQs/21VWWSoM2OqaS3ToixR1kDeq+MfbHBJlyWVCmMbvyucS6tKq1OE
hy5vYqvqY2kYVVlvHa4ASbw+TrE5HV+LBnNYXDp+29IyPkuEKS401o5qz5GJ0Fiwx0ekq3DFHEBD
TRLRcZ5KqgTmtX2G6BYGHnriXDQyMoqo2Uwu5w2t7fQhvuX0Ie9SXmqi4FU2BF5N/pdOncloS4yd
Z0ULEEe4nSfAbrLe3JwKw1uLtF0Jak9IL/MNx9MwNenrYuaXnjwtAGYxZgChXv3Yzi15R4IzwheH
g+EMBB+bIbP6Cwlc26pM+YV3dvg/r1p1/4nO9kopY3DzU7TvzYoiuozgq/0zI4Rv+F/GczBVHAVz
fknguLwu16ZZ9zqO4AyzHIiq6uFet2shtDssvCKg9TPS9MRAOuLtfENFTFigj5Ahj4GXCyLzLaCj
surbjiGwFNPkDrSb5GtsPxix2HwnKPzntD/t6HI7dfuUTj4zP1HJMMRR1SEr47P6lTvfTS7n7FDD
oAFxAjWi7++0biRD2QPTB+2enjuk+z0PdERQsREZtijn6h45Ki5qmAEI9TA7tmX0RBbYTpgszktQ
Llp9kxvu8fLf7X4jm9NDxP6Alt9RVjR4iUEluDNrSgxFxC4CTpg6hYTKxoAaRE7GHNWlpot+aoDq
2OxGB6D8lMcDAP84nvY6pPlh0+T1kNREKPoGnbtneduX97QN03545ijeB4o9cHMLYwlP1xB1phDD
Qk0owhpxPyze4jnrjKQox4O+Kp36EBjPrSVffp3p0umEZTY4g3tkDsgyVD063uGqr9QAM2wuGMld
oXRHg+Yt26rRN1IScpi4l0RQkOiFxpVNaUFmH+pD+jY9SJWuNkNRRQ1OsLvA2z0ykXt2xqLHpknO
f7rhYQl+mmpQFTvrj8wFn2E+porszvC9LZusYB2yf7qkeRdtuNJtWcOWTAlLEb2NbfcXJ3It5YAi
4P581A9VwwbmewCnkpGk0O/rA94kSnL0YshD/h7JccKilc9++f+e1SNfxzQAEzouIyBHHk4ZP2k9
Rh5Y6JMI6YoV9GhX5KGSnbKD9WfKRya0Yh6LK4lPyYKzgLOms0/7TH9xf2t+0TfA5/rnyeWKpV6K
g1CUBzFJcpgBZ5U06zcWkYsT1yHH+R5X3E2zKR+RnbGwZPd28ZhmDzobgAvFIzgZgRpACCr1DljE
aS39ArXo2YzGIDkrtm8ugiVrAEuWnWfRYC/ieiOp8vKJYMFWL3FWuPzOV5Zc8X5+WZmLQi9wLlJ3
jNOyqiq2xFUHWp5a4JDb5oylduCUPVe1wkB5KItYgWBsqELCedoYELhDNaPxrMmzsSfIxwBZcFSm
d6jqrhyd+83Ygn5/C2hWiU0xG3roA8B3lR3bFWtPxn+swo514qpHvDgbw+uVvNG9HKdfZZ4zc+yT
2lXZ28Hshx6qY9uxVVuoW1aSI6Kp3LNYwLoqrIw0u9iSEb+YfD7+IXtv6fLeWyyCD84mkZZjiXyr
A8dypXFAdYDonh+ZY5wnEXKdGp6LUHBOrtQP5LOpVs74zFfj70dAfmI1i6vziZyxdtDfNkD3vI6m
g+d92mJc2+Sg61qEtfcrg4Kxj2NS7lMmY4cZIQoWgsAng9vx6gzAgBmy4CcdKTyMgRGyPTkypszK
UtLAUR5KnmWovLp4q09ghp2VO0tULEINh6gfnimLX5FZbcOsh9Q1D2xbf6qc/v7vUlFISHaOI+uQ
eKH2xu2mYt0zW2R7aKehiFA4gm2Z2b1NMSe8cV+a/Dj93W14aXW6Tpdx8hQvtAN4PLaSg+NyCP1V
+8nEWCZlQbfqipyogB/GWdKjFk3tBjvkAJtTXnqzbZBxP0+tINXuoSkrYYXEOse4mdzxz5NTnQPI
TIWRYjPtkUxITEfyanl3kGmufsdSwCZUqM+lQkIB6KhAZSbE7PseE1mFgdLLyWNK33g08QQDsQ/4
TGqzdfv/4r+/q66ocJz59uB505oaIOOkFwrtMVlLBxSDNixatf2Db/S3r8l97vZmK9ofZmAHxM9g
eCRepTFuzcJmmHtBZg0jV68CEt2QdvFoAfoLESr++LT83xXNN/ntf0PAJJ5nChMBVBkPFkqWUrVk
LUFL36cWsd+bdcH2IOsfNBgaGJoje1JSjVjwJQkGO2Y8P0oCHmp28pOQIaOMMsNcs+ZiUYOE6lBZ
mmawDkBHo5PsQyY41M5j461v5DUZFgQI+epZyRUcFfnRwkRS9brs7mPPUXgMGjcFA70Oae/4SIHG
EGro/r0+W7oIUNHho4bLYLxaEm1DPdRm1omfKHentnSuPBUwdC3+1ofJwMFM6ZpUDeTNiJnNa6gT
Rd8PEc5Sn7LvYzajCNvAQuKXrwPjhTH9sEWAHrIzdv2F8tjfT1RyVn4VNNIiV9EN9y0UymSwHVsY
F04Q0MzLmy4C/v0QOqGnIzVQ/FqT+VNttqoZABhgEmGelAZGO+Lp7Zh2P5h4wznU7nkdD8o//7Dy
PREoRY2MjMBPnJnAAOtM/q77k91qmA/3KfeA0iwwRkLix7AMOsdFX0UKgWAAokiyoTIi8c7GVVGs
FARoL0DOxFhlAGWVVLoy0Nrj3g+8pFuMB36OyR5ussbrsSXWgtUhLCD8M9jhPObJFF00RS4rWHbp
1f0fpkpOnn5Nw7zwukMJAlc896QfHP2fxPo+3cbVgXqVt785kC/Mgte6O7kTPhO8YboSIbKjxrVT
QkORrxOlFUSrrVnSkP4CF55hcQ3uzRju0+IZiPJNd7AAHEe3PV7IRl1Okxty7ogXEqO69wSIEr85
Q/jHKpX8Y7dEjACgf7qkbkVtPFSf7TbLKqozhGzAyL8AWMfeLDNlEeOKemf1vKT7g4E6VLOgyzIy
5iBSIXj20ytxC/y0lAPFV937dmLKu5nAAmIj1QSD/14CsD0GkX/i4OEb4r3zk/RvXM59ZDFuhXyE
PdUB1AJ7mtUkp2omQ22Q23FmAaFEtDpYR4ivCAHReK6CcJJmIDZUOpeD+0GB33+cIxb8vxpZDXtw
vGgo0k65U4+7f7NLxX3254k/ecIHL5lI8hWZCY1vD4uVEhQp32aj13OfAgqH+hF1G7jXd7UQ3aiQ
4yByolOOaJBV0Vm1bGT5J/hsbbUI6YcxojY4pji+/x3B+BFr7uoT617Iy+ngUNg8mBnPniQsnutN
YK69qROoFxMXndlA1f1pzc59vAt8T49WSnMa5Mtf8yMuXE1cYpxDsPeFFScj3AvQZValFxWf70X2
W/rPsaUPT0fZObctyqAuzzdGZfOGvx4TWlEq6r5RaiK5qwfOWzwvGOyoorLW3FZwbKEt02aVU1iL
7Zix6m6Cl1sWHRGzLVsGIl5srY7bY9YFE8loOgZXyfW6VorN5F983ttITXFbDOz+4yqslxyPTuFj
xcjA6EmXWXrzqQbC/6Ep1LkpgivurCOovRDmRh+4WjT0gZZjKO9vf3oMZETGfSTWb/y95DDnWhG+
btLnlwRetYqqOuwJ+BIFLiEDQFveVAspT+Tk4YQVpUSplKVehmtAH/U1scBYW4cEA2pB+iMksn2/
Hgi9MA1UdNkTEIZNYTTHwjQoC397P0pztUm7wJKO988uRx5MYquB0cZX1rJepqU465wKEgvsjzgV
E82aJVHB234cNGw+C870BN8OWOiEfgfMjXmpslqvBWfIPu/IkObcnHwFW4Dl4qaakCK5EFATFOnU
qZ/tj0ip/ISApm/1kAXPzJFIyjxvUaeiwzrYtWtjIeFcVqqtDQnArPhPaUdOVsFuR0IsQl4YCcq3
8ZRMMs6aCjDZtflZLiAnfn08G1E5Vv2XgjoMArVc2+VTvE3LEVyNWudJmoSd4nMa8wPmfp7LJgVm
bfl2Gun1jgP/ho5dbm+yvbXa/ZCNl5t5IfKI/Gtsh3KTlmEQDroSqrOcmOlFBaNAxQkxgTFf/U5o
3OaIDrE1RSh0yudQ4ZcAqw2LxW31oburbkOmEy7iWIMRvY4H7bp3ig8LMxClRVb74yZO4y1or6OS
tQjilHtpVTUMEgEShXs3hhkS5ZS+3vV4y4K8JC2gLii6hdM9lsXQzrh3VB54Inv0/66v/PHSYNw8
4jR5lVIF9s1PCCZi6LG5qMbgMdTzSfongXASCpmrUGRdb/ROigyGOqwO3FI2kc2Sv6DAXW7ldkKi
iFf/irmFJ2KJKSxXr6cl81AD1OXT74kxWmr34p0530tDVpuaMROuk2qacuUQx/iECT6TDCLLOs47
kwOZ+YWQLd3SVzl2Gr2xWhOZzywDJZlRsopQvF++uOMYacjsuyzIyk+aFCHHDUx8P2k4iNzfuu4D
mOcUYvHC0veTlkyJYAy+CIXgnCpojN6hBWcPmb2Hvei1PRnRZDzTjrcg4GvhUmmKXmHjy3p+6L3/
SkPEfC6ncbXtnl4yhJM2DlsPUFpexp9nxl7f3oOHFx5JyRF8U8ItVKiZMA5DjKEHK09PUj/ApKOc
Y/VLpBIaVdw0k26cSbtSiEIFy5W32PT8DF+DU8a0h6eZJEEvLLI4v1bcq+CRtQ2a/PFk+jE7RppN
7M9fBqbXp/00/45XS800jx/9gj/7SAj6fZ/m35NheMI7M5YNLQzl3A8gNxSTwWaD7ZqegYFX2qn1
XbnOKmONLA4k+TFGnsho+4hzE01yqZR6sdSEIZfInhMKg49Gu3bzgt+cFt+M/CUZk8oUwDSOJq5n
2hHpxYa5p93u9kXmhFYNGVIPJvie/0e9sXeGLzLkuFOXUg2pQyldycBTdF61HSFTO5YANK+veHPt
W0BX6Q2ueV5rf5kXhHcCxslP9jEfQcCKnfcX2fdQu6foSS6bmWZr1bL4v62YrQ3SUeK7KUF4ABYB
zmqBRsEp61WhxkotRGz5EhTWMwn1Fh9/gWp6zN0dNd8Psw72JOfvlYdem6Z8fwHVd3zr4On733mk
Px4QfEzUQClxIcCG/Jm84vFw7mlNle/+x5TeNJ1t0fBEnnKA/5m+Z+Sv8BEFf1wNwwGubDXXGNj5
QXQvvdHoviGiuzgDUySQtvEMXUcV974Z0e42kxtdPXA3ebOQTZqlqqVpup3HvlPO7WSX1A7flvQH
AVk63zGgm//5N+rauXohZVKlPuoAf0vkgnJbb+Nfc1ekSKWOV00yWx1PKBrsh9QAHWm3kcSIQ/CY
aJLbuvweCzF/ATal5ogQtaMQ5N/tPXRHDK+SgH+kaH4zswHnJDVXIFunERU05kyBVeVkqBHKaJoK
eCtbRnfy+b6KExSUxH6MgQC64AcFvTj4Twe7xiaodYKPM71t7yKccQgNmB+0ThQUnSVWXcvccvb7
GH1/JLG2U7Jiq/GZcn2K4I7NtIlYalUDTSANi8tP6gy3HxYNLi9+CsJqoi7aNZZtcj+P30+lpfqa
QeugPd0VS+HjI1GZ229mQe0W5LqD3ttrvuWgrkd2lwTxgYgynNrZQ3INmitt3ZCEkFcorlF8aOVr
xwvI1E6r74x6E919fWSQMgRjHyDt+ZYViqgAniS4bIE62yfcvuRVyZki4+AwsZkwhVPOCYLEJVKw
VsJudffLeWLwC7rp6A+Ivk/uC739Wc13JPDMP5ZXoVwdD0iggogZj14cfiwoM3xca1MHH2LXqcPl
zPT1+uBb3bBlesVHafL1VfEclU/lMzaq1qGjnp3RjpLFlK+YnbJ0Q7DUUeGuJd4D8SMK7uSkJcjO
FFYjTlpaFNnKZ8ViUR8Z/fmoTWaXFNLPoqyOmBiMfjnQeBJxzvk7FDdgd3HShLCEiQLzE+fjQoCx
A/kSe98SFda/mwPU3kaSegLKrJlydE6iQetfpgH0HRijciXbFYfqqgrlbS2q8B8PiFiEKpFjMaj2
mYylP9NPtQjfunIBrlfLt3FiXNlrR6moGDzgDe4nBqJ2uCBNSM2NlD6SjQad/kOX0whqrmkWC5QT
8N8VnQRm7ywoy6kHc0hZ4LFGNvBnf03oUPonHyP8U2x7ActybwnPuiXfWi8aXk1PtZKxZfMlGtk2
rQNijKHHGQKBHcLU4sVQBAlKuc+g5fOyI1AmjwyeYGhR3ee7lnXtetIlatWrKNI5porTgew8DeCS
MFvYbpLvghfFndWdnUB+HI2FVXMl7EcQIaYehyDQsKOnd7DVYfdRsm+C1M6j59ncXRcNkxnffL7P
fsV3H8An/rd8ypbLprdA19odrnKBA8BqhcajiFMq/S1PKj3oUZhZQvrZBhsY1vUje2qrHQ7wfVxr
HMo5zIq04T1tL44l0jSPx6BhzR0CY/iYU/pqowfIxy9T8LIycBVdt4Dhor4j1n6IyEFX/5tBcgps
PiU89SA+8eM34Cq3oF8VHF8+vrj6M0/cMTWv88KCgXqtnKUOfAHhKnDe8vRFFLpuPn0tkX5Obi1i
2v3yZiPD3vCOZcbpaf5vEwqXb30wbjOfVxMSRgZIcCY+DhAgyiz1Vcumq3OJhkHFmNMwvRqTi2tW
T94aWkuLbYhyQzdMtPqs1JeZRayQM1YsyDpXcsOCd1+vIELHW73NF89i6E/F+39JYfbOpybavtqo
aa/1JaX3k/F4fO3UjP7U4aH1Ye7EQ4B1pdlP6BKFbJFwGPNAC8Tz07wbsWOF6IRXUbv3p1JpyaKd
n+qnXbNq7eTIqUROmyX3Xh84ovIW4nopGXE22iCe5z549V/rEkJy3IKNKYmGIyw+/oYLoY66ZHyO
kkxCRWMOUrcI6pFb9TRB5dct5KYbbhJODDQplsGud2csderTLyONMgbWZdabvQ+fBX/KCKJyYaFf
916H2Bm+kliBDQv5mJI7vLEZcJMWD+mz3NmbHr1omOSagYw3H25Y7PbfwfFjK1qaE0PXMpr/qjBP
an5PbzQY1Y1uq/IV5vnWcDYbZsCEsct8cgiNgtz7lkNWquYz9LNZdcqWUl9rbedU1nbl/H9UMCG3
o43pNXC3/J+zyHTxfu87UWPL884BfQE0yMACloeuTkJYAXcHm+OsYmO8GWVKa4a19H2fn60C9W24
ueEsAXPqO9g8si4p9L4x4jNiWuCzpkAxRYWcZCO5awS0j9G9aZwFK0RPtB+jSysxW4dy+YY3SlGN
2lZwol5EFz1x8NSNEGXafkuygSgKP4MBQby/1zJWtMq0uHmA3fl7HG3Tzea1l37tYjwvGdE7V9qF
e9yMLrhamefFGhFRuSKmDWelGcB0bMXiDKK3X9C1Srr+KFlwYj1/0ErM2P62aOYNQA4CCpS+80bK
FN4DElp+qLk6Vu7i/aZpOj5r2suJhNVqecccPiM0gDQJngbEflo6/9Ii67YyMyZRm/5SGM3r1bxK
xS6j4C4lTOCz4PR55/4JXtSEosTQAK3Y5oRiIlxFtGzUvtYhVcFeHOsMB/PUflhaXprBJtQn62bH
ZG4eCKCIMKJEU8CbO5BuIyd91+bc7WY9ZLUn+PzL0uM675KjmOvYsYtxW/iX3xZIMavO1L+Vtvrg
xoF5DblKWg5j80cv7vmhUUbuAd3D9Y1ZdJ0lcBl5j61JQnqpBGrDk/AK8985TQr26S5iE4AVLTa5
zGwALGt1r4TnDr0U2ezmyf+aWfXWJsosDt7h3wduLLpN4wdQNiKMab8UusLksirkzXgcRHntn3+2
W3CVr+nmMLWB0PxeCAu74D7iwY+Ez+TtqYM666yAdR60HekRxH+8yDP1EDZeK6dVYtg88yMMeBA0
MVufLYZBYX71ibrI3cdddt9lYxCWNU2U8jdY9mMt6aG8bHukNV0cUB5H2tJ9tW6c9ATyGVN+AcCe
c+nbnnPaS5FFZ7+UI+fam8RHScaT8vBui/7D3+zHHY6NsDb2y7XuDKkxD4vMOwdkTY+xXJubfbBK
8q1fG+EoIs17Qva6zqJB/dClFc+rdNIGxHTs5uI4giQf0jaOG1X+6RXcjg7OhtBiDgdqztJjrhMk
LzlL0JaEvw4Gg/dQbqbHHixW+oOiFCZMqyWBkxS0hyTSSBcAEVzuYuL4h8wNjyNF1gOWgLBaGrDb
MA+noyJG84NMvBM6kUe37qTdUsjwPcCXD84y2Mh/T9fFRQkmes6ZuL5aQFBlPMd5/+r3uFONJNB2
sxzlR9Bb8l5dM9fHZnMbji/p4yu+t/XH46VmulLOfLJF8muDRH2UFx4O0Mgxj2sKZ5d/tWjT7WaO
I1CdD+jnRfoRa3Q0NB7TFuOJOHR42/pEsI9jpPzzAzWc0PN5VzySaHNNWydSiUp/86f5UanlipsQ
IqsHt/TUh6k//JQO+tkPGUoZdD2uAyHJyOShCPNsS5sD71K97L3LSopcilQdRnv4QdMf75duhMcG
V8hKqqHWy7FjICh3N0652cyg1N0DJZ2Dvwk/sC3ZuCtBSkXlP3s2jmUN2r3feMHLM1KJLWkoqE8x
dXEfHbTcWPrtdVhOLE7y/21Xf/NY0Cj0lCOQwsSVTzcqmbCJRIKu4RKlOpBiA9PAmXnkjx2zJlNb
gkcYKNhd5q+ZU/+NDE5MfZ1VrKB3YcLV1jUmX92T0f1YILMNxOw46J/T5xXsZVUgjYF+FWGyFpk6
Gls424dQsotWbe+Wd/GnqGZGESLDNhp+naZYpFbGD6iQITY8MIvYGrr1J5g/EUivMq/32wj9+JVA
PFIkwV20zU57NF9u0jlYp4iHHEuIuzMZM93/6IDtWYWRCKPan6kQ0PGH3iiNGJK7c7URk+wAMYEJ
QwzpHKlHIHbBz3NSftY9lYePEwA+ivBjChBn242G7mkrfjHXKkPJyXHrS96Nu7KzX8zj0+oC6v3E
8DMCSKEK/t+Kz7XOPeg3n5n7I+tiD2gz0WgFot6WX04H1DL/Bd2bFCoUukD2XX2i0DsqXYYXhIiI
+V4lB/zFLOv6dKK75tj18AyvMHxDZSlCtniVFxH6nw8Tk0e9FUMVLUQsCQV3FZRN4RE+wq+EIv+1
jIt17hcAz42wz19dsPXUZ68ar8ds2a+Ys0o5mRUB/trQyMcPjYZh4nvsAfH0r+fRdRswoHxnTw0G
fmG8ICBBgNoJE4skaojENYEhuOBOgwQ3N3VYFvwK7O6sIOeLFif+rn1FUkuZopIbLgGoQyTR5wVq
oQbyoH22YoQCgqXvWnJSvKrlapZuhlJY+exULJZcZutrQ2g2TQBOSnPBJf2aWKvyhvhlK5Bu2jZD
70eVEaLk47BTqkBrB5OgZWmTg0sLiQmRZWHweqTVWRiWKOe0guYYw4Dmmr0fB2DukCJDDLIjHIvq
SJfdcs/1UHonO+4UMX2tiCDDBkKIeQ0A2T5ELQy50l6txqj6SGAsqDcJjxY98yFPA1AedcXGkVz/
CJm9UM+IHB9VATO901oaLP/RJulMibMON/iEyIDjphFWEnz57B4zmu2qkLHpWjTSVspiVYGkGTRz
/86hxvqqfwhM9gv7U3lJ2wFvxl+ppCNbSf32piTpioIS7dEeDgnO/gmgB16dXMjXt0tx+EqViMno
rKcAPVPIQeYrJOTXzTvYGl2ayxGvBhPaWbm2xm9HKfG+0+V/ALy5x6ao8yLnWAjnKQKKfpPKPBUG
TAg8akSP8FlyvyArg6AeunTYybyEAz1kixf/BJtvAhDC6HUSuh55ODkxFjRG+gtXaHvAZXf0SuIQ
Gr4RQ3PoqgbX/+T+1p5FSXrzX6pOx8c+zGE1x5GnmXCOAnq3EZ43GaqzZb6YLDEgOwuegFj64VJc
gbHvgt6BLqNi6Zk0aNttf8eY0e1J13qh+1S+lROxE2s93RvvoNF2Cu4iDhT3enVte0uPT0gvHUt7
6Abkl+Zs7tcULROjJp7PsgOozKl9xlfnE21xp1NPdLawOClQctRlErKji9NIgND/N3bHUQIeoT7D
8iU9D1slGJ+4deV0fe/V2dySrpihDunmf+rWE/YdnxZGkuCdSLTDdvE5cCruL9/dvJRKUGNY8Ja5
sK03wETEE1k7O4TZre6HDEEqx3elWozoJiy3sYm9aSxWXP+7r/SY8SenE6Gv57Nnr7nIKDECsYAz
+uRGgUfTJ62K0V+HjQ1Ds1l3Bdg+oaNpn8ruyBjxLxAJ5HaS4hCvuFGY/QY2oOdpzq7QkruwtYwR
YRjamAVqobbyabd7IfwOCA/TD2CFChZOEZtoLwL0nzcfqymriud4PH/YHMPsPjjJeEqoa6fFhHry
Wbw6jMHSxRaO0gDw0PD5sxzXSwOHfWH/3RpWZxq09hCrOEszRNVgNkGVw3hbz19NxdKb+meCjJ6n
Dv31N18e7Y0hLBl9EUDh5iJsU3dg4FUZ2x6/fnZxYsAIROPtxqvLCzMn1pweQcfIclLrb1Ni/8HN
rnQywKf4GFhWnLEh9IWegG/go6WOsMbxFMEVq7AKCC0XnL7q9EkLXEMIWqrvSCeJsiPiDIz6deWi
ZWuac8EfVRkHlPq+MsM9BxF/Q5HApQwMOwez0hK9McKWauNFi+eSDsldQqlGf0eIMXIBIJ9ROscw
PsPiY6R8K4MY9Jy8QTYJVTaICzsWpyIQvvW6Tz69I1aOx2D9Ibjid8LJd1SBsxu2tE7gMCs8CBHE
/NzGi80wkC7sabR6DpweuS0/6Ou9anWhVXsxu/FOLkRH45iPkPOJYL+5r3ZK3ioC2VfX0sOgcALc
ATA/FpGln2eouQUgGOLpnWg0JQGI0QJRmrRD3ktEetiRV+72FCvdpMq0XiFJQydWf4r6upoP/WEz
f0MiWm0BT9Qyia6LsgtR49ksDZeygLjYtAcWX8DPS7t5LgO7tyFxiejSWugKHwL75K3orNhRWD2u
zmcvQFwpk4V+CReTjEZyImVdyUc1e3H3mov8pWeU64ISm9p8D7YGIbROiGsH6ZJsd1aK1KLIdgHH
o5ZrMJhfBt2YlukPPCROhx70zvwoyA17jrSBOmIuwfrUIaWuoScJoBpRKEtqvJjXFihXuMcpxvCV
iYR/+QX+YdxlnRwRZtAdT8ot5uNCqEGL2/afK1UinVSVU+GEE9kMUXlnbzHAndTutPpd8Mfabh2R
Tiiw9Au9em6aRKxn3usnxk4+QnhbvMbTdHebYa/SP2lrfmuOpEfFjvCKche/pb484qW0tHmLrEQ/
gasSuMqk/IAEnyOKUf1cNsOPqd/hVyjbvL+aU4kc6P5Nh4b2LM7Npvuc9Bvz3BX4rTBomt6n93kg
kXieGqSLxDcHzQNQtfVyHM4RCrmTb8W+Pp5+rO62DF2qkbYjupuBdeJmlFi4KwoJZ5hK5b4OfbSd
5R4amcba/ikOGcyHm2NMSK8auSjgJ8NYExLRGdYhgZPTbCn5QcDuPksUUP4WZprZwvE5gwfMm60g
gV9xsr35kzDCugKprp9PzeH+mTaDEpQ9LZL6clUvmp8PM+c5i/JimN/OQVk9cA5mcyOlZiboT4Gl
SmASWUqtnOQnfVSkZvAsX3dWu7WzpmEHe6D6poGq75VDJE1/VyoFlPoknC42yxuJEGjbEWCNDAF6
3y0KCr6XtgNoUi/KjIjVNO4g1jj4PN0njV5+HpTJ72OS9a1alQsYiWH3oER4fVxqyslMR+DcBLod
ux1/1/XSYTp8WKi0O6EJdl4YeStSYNkeiNXqnV3+j/hfV6AtY2rEhqQvB6PO6fCvLRxly4h6fCEm
LSXwrKmWuCtrispBLrqiBBnutmN/LnzNm3TGvVoDtnbHZ6hk3Erv8GdtnJWNU7iluN5/iSnD1VNe
wvmmydTf2PyA1d5O5gl4592qoHUHNBtORlNSOTj5+gJyz6cmF6s6Fvr8Y+kTrk93gk7QqTnqC4VW
jeJgLNMPhnnbRfrrPrUhuJ6fUuZq5UMaeoooj43k2UuH9sNA7eys8m21FpjH+FyHrs2PBj8gjsMG
dazta/hTaDU0BGLf4y7tkv9Lj3W1jjpjNIBGRRSjf93Ev2NEeY1hDjAYRZPgnINWUt4KuD3j9HJc
+awjn2+XFWd9+/pNnHrlhHMoALLE7r0jHskNT9wdXSDEVRtVlNgdaYl7ByM86EtQtgt7uScsk9gA
WexHqFHwtoqSssvK+6C0ynzkbT9K2neORm0Kfqhw2+iLZayvA7bmdxW/joSXha9huc+2gWdNwNyb
xarYd3Ucs9Ll8RDMWfTN0wQyEjW+JlaNTsVf3Q8DnCJoZj3N5chYfojBmjratXXxnRq7f8UC+my2
MjCTfKpMzEgUKxhPEHlXcsLB2wBTBO3gGRPVTxqEygqIEWUhSNMEzLcTvmkuaguIkHlsx+HarUmY
qFMhamp4U6z+U6WCSpPK3wyydyGbBXxFlXN0tZr0BgLbMhZN7BOeYrR9WLKCKqD+SE6LzKaPFVgm
zCsfC+y723nEZoIfK4aaKFeVBuEccvMLoOJEYFIVzlmiNJmsohg88gdzsUXuEnvi0ha5ThJd48LY
WQJVMzrXmPLdWpfednr2YK0bpEnokG7DzVrMXeHR2iABLRvF6rvbjdGeZcOx0p6bNZzv7p5G3WG7
C5/zPMAICONsRGhII9o+r/d6q88vxpafz5l9RIo3UvCEkwN21AX/jAn1OVPgdrlX/4KT2UoWXHYg
z6sNsYEs8kuShPtNH7pvB718p0K7BcaCuU+MendDXC9amX9V6yGnb/CKUcc92qYg+rLQ3ou3p5IU
u4chHNxWuABM4FADUPu9DBnVpeiGBGAhNY7qjCtmULRJKQlKtZfCEg5B5GOIDVks2LzPYTdaU27M
nJK+Oi6ECdZrF8x913jMCCr+tSAjN068DSizY+PuBZXkwKT9ukx45f06RGGS27h/ou9+0CrMumGb
NK/2CkrAY8HzaCsctfqYTa2zLorYBZ/lZDKQHnpocq7reIv37cUZ2AKd6SOgF3OQHgexu4z+noKi
Z7/qJ8glv5yti3IvhQ+2er7gSxcdBGshuwh0GpWHjrVwTmD3wuWTQ0TDv+3p9awXujZijyQ7AeT1
SoQmzdLcuMNSYNYnJEiFgxNIaWUuO+thBX0zLiXTn+2ratDO+zezGhjzRAJeWLuKDBERqHsEFVN2
LwussXfG1MRPyCCUjFn1VkP/xKFQAmC3ppieKiZ/zIHPAPuAurfPNCTXLtKCanRovZkk7H50NqJJ
nAj+8S32Asn46z/f9C1P7Kl/XfL+x2Ne2W2zRgY9ibNg6evcAkcOVRq5ZdF1lCpS+2wnfbg6AQKd
Nc8Atv1+cIi0BU95BV/cZ6mvpq/BjdpIds7dFJa58+71hgmdXNpNBzpeLFXbh6sK9tEKb26Ee/OT
EAHHjSh5DvHPDxa6q+e+FwHBNajtyumHyu8MFPIr6ofafC0bI0PRBprhnLndtBD7JexzAVB0Mitf
Ul2tNWKGgi+rJNp0PEVp9uG7XqegMQoqCFZyTUIxaMHnHKY4FTerGI4gMqOAuHYcQB1Pndtzwa68
f9q2oiICanqEz2VMWFi5eT9iquLnJgsh49xiP8JBjcfktU8Xee/9BGIAj8gGKB0kNoHFgB8EzcDc
vPOI9Q0/3JjinouMUrNLiWvDimO9H/UmB8IvjFGrTgo68wJ2yvNOemZx7i+r/BnQAEtoa0/lAcDP
HFCNzd0HlyJQn2CWdQbHrG4+m8oXaMHkTSMI/u4JD4ARDRRfYLTVhYsAxLWg1pxkW6ecNoQuQBgT
RCDfh3kIhYaUdEHz5RiP8M/hScCbpZgIwJfuCxo7Ekr6suCzN40uhtxCoaaj31WntN2SLHyPMU+X
BuEVwigJ6yj8sTqTMd+RZgOfA20mP4+6p2/Ym8MNv+0sylSxWzLqqwVcDa4FpCc6tKu/I6dGWntB
LBKxO6tgG9tmdtiIoHPbIWJ6s/3ZxmBzj9qXirOGsDhyPtMT/OBkmufnAQ3Rn2gRfLAyXJR6+Pai
LP0N/4HlvrJJErXk8bt3grDt2E0whFKnale9QNc3Tn0vNSpHzxee2YCrjXWcs2snkrWwpBx6Gihi
3u3IG7qfKz7EGZmNcGP6z4veW7Kpe3LRRjV5Om3Uu6drMUdQEh0yRnzHQhHSlPMoPjobv9Y2OMCf
Z5yaLKRSwI6xZ/GwSMK8Mxwnv4tNplNRelm/q0UkO/LCFwVlpzUXW4ga2bGh1O/a309HYabIqX3P
sdVCoQ+f3Lxv3V8qLYGHAltZbBehXdj9DoPMR2WdnLY9r1yrTzpptVR/AQyTBPFPQ5S3C5HXK6PE
o1OzOPFWcf79k23dGBbFKQw3kikfl0nFB/kWUnTM0pn3ZFFo/b6b5sdUyteGIqviHZPO6770H7H1
1nOQNUZyGypsfpMM5lZmbeCw7ne4jb3YeyltL/kQP9yDOGPQB8hozZNnXlwO54VUJLvTrBjN9bIr
zua3A3ZzxBFfQsyLpYEoI/XpmlD1wP8IUg/bgm7ESKFaSxjqmgu1ZQfwwajd867foq6qWC6DDbna
8HND2q3CguvYeyhyYZwAT1O6inhjV/nfeIjCN5c2Nos2NYcnh0knc90GPZSv3hs0g+Ub4bgc2FTq
4b9y+eUqnMKWim0LklgMU7XX6Lg/33NnWJmtGaOLr4HfIiA7UxplgFmxAVWiimzxfLW+KBgd0hLV
G+Q5FeDIpuYM3iEfbq05B4BQP+ANYz+tnX4eaw/m8UEsG4dZbPa86NUfczdHFUDvqndKpLgtOyRd
CF2oNZunCukSqCYDK3zFcagIDW2aKSH2GWVpPs14i2dbLlaEIWNGYQk8hJfmmppbYPauITXUejh/
cWWgucswyaJLeGnwDR+r9NL2liV5C1wd3Z6iAmQJ//CnyEC5lFmubVGbCexhk3S5Pptn8S1j+gHt
FKjbaLjtN12sxgioS2NdKfnTPyM1/4CN/BvNhb2r0FO8MMWcTrvDqjeAS8Yc9UyDSH0rw6Hn/Qh4
HT5vmns9qqzIkx8A0M7ourR0q+TJdpT8tHDJnQBzHHRbRdbeLiu9RkI7rJY9JLezd8fEHpT/mmpL
1R0BRWLrSNERhI7j6FtVSlQwjBkpye+2u4yzHHOzzjHKJFdqmDaDGwXuDXLTxPGR88M3qR+aiwCX
Up5vmgj87VtNkkUK5FYtoOrAUx/nrywIr7pBkvbgrzQFflpKwlvmcNImk6UdDvTDHRNpnMvdL5qZ
R3zl1vSa21410wvrpHfAR6F3cVM/STUQ+MBjGe0fPd5m386O6rGnp/oVdhqnOaQIKsogwQibFHgK
8gJWnGQ0N4vq9/pbz4CPZ7vBPVoPkDwNgVkSq3UxxygV+FJlSv36ePLw8EL4a26IQ6evVUw+fMhG
r7jpk0bbV3IfJbSwmN6VRbQ676v2Iju6hZvWmCKevnSIhlIqqW/3DQnUDW0WCz5S5JajoVIbRbda
OOD/7cFEcC4PTqlbdcFbOONo55fZ9QOT1lo0hD8J/iXTtVFY8dx4jUE4G77Kfgirx6nNS9JCHFJE
7oPet9W5aErVVAUwQUfL/w4NEtQNF3M24qX5mP6ccpmsyIvs6DTXaoTODy/JVFU2PQmaoOD4+neX
FaaLn1sKTM2736MigdSGUWug0bd3B+7G93H3stfT/VspxznTVcqNQT52sftoI+geRKjf6urZQzZ6
zttEIlJ1c3REikwlIp3f/vAnvY0ND0rYeiHEpwjTWpXQ3qwaZJ7MMLAFxT/y5JXtoS+UB62bHlfh
u01fLDIMMo40XrdS8dOXa1Mr65w6icfJ0cwTIkBjYEbnfhCDPS/plbZxpYfZ0+0H7/wfbRR78LwH
htsRrzmhHPzwWz8MExC4Ej8DcALkwBjOEG2rBwO1TpGhFcdzw/SoUe6BZmb5wyq94bR5CtjA6hVI
bN3Aw51uyyd4gDZJNfKQ1tYTjchlUoDF5zu/tRXVIv7QdWfCld5iqAU30Ko7ktMndbx0srkvSomy
KDnVdtKGrbRisNGWe6hrGVFEjtPuoT0C8xQgwOG0bNoNGG46zbtIogB806LhUugJsCO++Rvwl5Bc
/TvOxFJD+aiu+bsDCqVrwQNh2a4/yJkOYzmjOlo1XnnzNskYe9b7R2V0fEWfZubBwetTSN/nbfe3
GADWTNl+ZZysHtxd553IyA9WfudkTpUEHWLmQ12OwUjKnezO+K6xTwwBykhdHbUuxLgKP9YjsDiP
BBFqRa5cFE7g/xcvbTHZA3kY/1FcPnoTX06pSYUdunOh2YhSjUdU0HQ9iLNllZAN5rWGrDVFlapD
SxSPXyKR68OhTmEVa/HdSJKimd/S157cTI4yNbQ7WZAdSoJE60dPlJLL1XeqnCAkLS/fMf/JV8p0
rar5Zdd9kQkVv/x/Yo66QrG9687x6tw5V8ezv3dYtG9lxxbyvr+D/PSDxjqIqM4lC0B3qVHiJiEm
2UgGC40NELUBva3iN4EogC/Nvz48+Hs2GcVBcaHfR5Air5I0OUCEqareXg8zqo8WtPrlk6xfTrLe
g3Qbc1z9Dwt2/63ZxCKgvVVdU86fsCFvXfsR8Vfpu0jxeTB0bv3U76fHDgLze2+qCUNah0xhJ+6j
XTS5g9eUthcxa4NiwDw2oPG7kbBgLZh4WeTQMVPaGFhxe8h7e+Rp4s0cBKhft/hkw3HfbsmSm3VB
x0OIoHYWNFmrNr04flL+zeXrup7mvw2wLnmIktPc0e6Mk44gQtfV9Ot823wlGc6dXsy3sHEflM4d
xp1SOZlBCABHCtrytHs3Cix17RS7XsHfy2rT90Cxj7g7CNC3Wp/wFwYKb3vCkkHfD0zxgGd5LcLf
1kbTOVu2L5RxKpbPj6pb6YeV0kQfkI3Rtvk0DbK1UYny0nLcMXPAkfF9vwOkbEctVf8FFn13gTci
FLKKK+BuKgRT2ClEAqRKlWndhYeWD+sZrKQKPnQask6+xps9I/BIhxhgi31RWNaK0nmtwogTYj8u
QhWgPaVxAU5cdHTK4JbUxN4CLnDx1PpWM7DzZwWLpbRfB7qAgf7WUwXp+N9QyAdxObLtV6wXD/h3
YuP/Y0/+b5RAN8ErNp0upz+5R6oZlzLXVB8XgpFTzMgfa/fXeaBMiG/QUtDir/G20uAkNX2ZxK3I
Dx0DBtRVB0zwSO4/eDN7s3GLuXph0x0MG4L8OAexrG0TPeht3Om7xO/UPP1BfUwTb1l4uA6hAkkC
XiNDAYu7mXSpb+lWN66WSWaEm4uoYZTXiqwgRDmsVhsCRIglFbUrG0/ZKndU7jeeof+PuspGy7I5
wh8y/b0jd1z2kgvTwqEN4YB1OwZBsF2euVxtWSgBJz2p0+Jo725CgEmd8+vuONeiJWfrfZ4njIrP
htQGxS/4n+oI9R2X9yWXYUR9vlFfG3h9cS3tE5A5uNJGZDk7s0FQjygoIVDd9+bofx+0/nUW6DdE
I7fQBhoJm9ZDzfMsrQ2mdCnvYggNZ0meAWJP/CG9buV+TYBeeEdYoX3vilhcQzH5zHtBdw6oc6pe
g6FYuyBFM7zfezB++2qWznhGlNMSvqKOwyLpWY0tkUiXqaEFc1TwkkaniQGn85o7kHMYi8/iQQgt
rjUchLtyxeaO9KXFLYXBCWk1qWJnCkzaSmwOCMN/8yVc0FaOWtEcQ4By5eRybYCTJ+O2iDgLloPM
BiQ/tTjtPHJWE23WsLFyv/ZhJqAzj+oAUCPvB+L2XASp+1pgJvV49gzBPblSlfLC/euNhgvi1eqO
bo1oGwDoBB+MsNzmlMAEkAdSVZTfTOo4hNv8lVk4xK9NE4rbULkheYYZB04PUDVEodwaKjAtirgJ
qoFfzn6A+n6TngHF2gy47q+BPTNTpkgtyzAU4dH5TyHlYDXHnpfQrDdXtyth10v6kcMSsKcJopmF
5vIvGCsVGuvPKOsEEHfAEgmPniIoMcdggTo9IILrtnIw7VdXrsnDsnVfLDXJr5r2V+rjjlJd36CO
tjhgMjORieDhiDw34I6ZcKmIq7opPyfbQPxLsZ7i6mWFIR6iXDyLEHDmZ/2dmATiY+AtyrHI4rFH
2hsQjF8klUMtU+Q5Fq6ZB8gLIv3oVLmdNIWyENeUmR3h9w2GRFUeXdZHv7WLOUjbf3i1QBhWhoji
BR9ssF2hdDjV6deYKH9vKF90f5xiwa44Y6sT4Jm7lY/oUZqWXhMKLtb22/OYq1badfohevs4EThV
i8SC2mS6aP8Z0zAptsxU5BXi8TRk+WRT7B75r2f1w8O+4vb5U4x1oDfy8/EnJkleukMICBgaquU8
meQxjSFog18NJTT5tF3+xeoHTWaSRT/h0GBm6u8wgL//dEADOswDkPAZa852WWxcO1VJM7zbYPvi
gY3M/Ia/+nV+IvCGunqr2selq20DEsXAu8C7KBnxAQqK/3m5NCvhfQMGCMn3MeD4vdnGqRYm9Qsy
km4Qr9ryA5CzZ3t1kNb16ka1s/9bk2SUWWCWeqTJSvrBbzfph12dxUhJDkz7YWHPNp1lbPFAOHu+
IKLhVpGhk+rXWg6RCLVZVJZJ26LgARz7WvpKfq1CsjIcOgyI30CVtxHYzo0tgdHvj1h0x29GnfEa
Q1tu9q5WiQ7Fr/oxELVG+gtxRGHLbTxK3yfbY+RE/c39unYHqvoPA5NzmqGt4++RGMKTqKN1Dpbz
cIY85iiUlD6ux+7TfiYOwo2kcf+nAQIb5YTL8oTLqLFzViGpshNRthyNiO8tMZphXZqrn+lO3Hwy
c2hjYNEHKRDrKceZOxZZwptgEJx4chUPx1LowKUHrhrVlER//438OYD5XGIPpJEOHUIkT7RPQhi0
UXgyWXSBSDqiRm3ioRwdY0B69PO5O40Qi2E/m0LO3QuLzQMW+zuQ1H7/FaXUaXuI9mEHnS/EhT9P
oeLuS1122fUzzOEuZPW7Z6XPve6wsmmHwwy/2sSw5hk1IjeyZTz8JCs7NFwEVWsWVdbukHg8i3Qd
WbM9wdk8IEH75OzlfH09k+fMIjEt66ITZPXBL1wNvKSU3OoAnbmi0PpGifzk/VJq//lMdVjZbamd
//QDENeXK49ZmxPAkOYnMziREp1pQxnKTeIc+1E9DyRpMKteZnOa2athWkTwQafFZDoJhVnj4gfa
2JWBX78U50wuFyvv9DNms9geQxRJoTbkLS9NlfqbK5gOSTCd5QOoarOH7EBVIMOlchcOZlWI4Irx
Flw7O5fdmlJ20dZxULDxGKBmoEDuoz86LyYX3H+V5tJ6hkG4DFDB0e4Phi7DXalUWJnaXdjwyRLk
fXwKiyHyMay88nFuzoHh8hoZ+hj0Y18BeOS+06fFuP5/MxQxh41OpBoRgXyk3PDqOyV40qS5vXna
CoJQ4MawA/dAopwVHSBLCV02q1JEG6qLntMmio+JGfsIg+YCisOu4rs9/Y4jni/S7/Qbk/kvrSWq
ZNHA6cW4+/bpo9jeitbgTX5ZD1bWnlEPNuhHWJ/kcifenu7rwQ8kZKiXn9Z6TP2SYKV4md3JVxce
tWTria1Rg5ahhuCZM5lC9hQpQfjuhHEZnQYR97NZiVNSl5dhIUNSWkzwLCk5nZwA/bQtDnpi9Ac9
UynbaA6tSgsscislHH2Nakh6l5n7eVcwkfdWGIHkC6bXOM63tw6qUNewT0yp9oHjD/SHVXODU9p0
loxDJmxyUjYhbBjCGpW/BsIiQCBlQl9th2wGb1DnS7SJPZ6Xp591L5mlsfNJBo2fZFJEnmTarIHh
q3TBFTzrpR/k5Uexg6pAeFDe7FKaKspffpaQoqgeAmzwjvCo+HiZQoUpqigfYAy8XYeEkrnUolJ3
zND+EoANKF4+fk43HC789Y0owCFbm/ipqS3r5LCEVs0wGDB3CNif6iP2uuY4k9SHpKMEpEwECLoL
oQvlMC4u2Z4C117vFg2AHPnuBasMvUVpKFYsPDvEpCAi91h8yu0MSD/7I8Yr2DCsPno/kd3aBZbq
t6BPV8UMNOjA/LrO5+IEXVSC3dYDGyVQYoQYX9e78FJ+muUj/rVzqegYYd59h7zhK2ONBSz150au
OPJ1rKr0uO21nFuZR8LqZWQynWXadg2WXuqjQDxWVhb99nqXpVEQ4Tf+GGJMRt/T0zg1pFpTFXus
aCsE39aTKW/ngFKkV/EuBmuN/g9riPQfid4eg2p1j2yzCGtJNKkcRfemq9EwJ61T2TCmzuqW6vgM
BXbcC+C7rPpf23R3jfSVDYxlI3NKvN1zqLTLtARH1hB+NFs4vND/eeit0WbqSd8DvHMkrLppbFfw
DZPzfKbUk6Tocz+sgqpBd5vujdQ5WQvPkA6lrSctQrDuaejABTPW+DhI85DqiTbuVDd1lNpN4Z7U
6eZkEdKwyBDCzz+/1MbN7Kega9H6oEfQxb9qkSoR0u3Mdguo+uGZBQwPOlbZSuhdC4CzfAcOU48w
/8g8T433kh4MV1gFfpZAV5PfB82Zj4J+IQ0RX7+crxP19iSGc6f2vmp3WptHmZdm8QRR1Sphx8og
6KB9ET67aECeLj+9WXsa4tJ0zFLqesnvOljag/JQf7yISKFF/QvwbbBJZOhiZD24xMEF+z1iT/uB
uA0hSdPd3jHp+fxo326HG0MpyF+vmd2C5emiht54GZXPu8WOQlAAOPo5LjsRqEwhm0ve0KioUpm+
6FKo0IfI/GU2UNg/JFhM/qem/LpTVcMAFYVKDi2vdCjp2IwZfm7ols16H5z9oqkxFRopDnj/NNZe
krNQIzHbukQesSYvm1VoMq/pp/PblOMkyv6oT3ZvKH5VfmMYsYzT4DLRkiE0fbyec91bgtOM7gT7
gxSjYLtE5DO3lqxedB8BwtvKeahIlbpdjehO7t6nmegq3LzHBZoBvRAE+uv8RRoBAg9mxHBvfKzU
TSh1jGPE4xj3HPZ1EIUuNKPdZ3UTZfSjnw/eAGR1lnzRCrrIIkCVvpoT9fn+mHhCLxSno5bnAZy/
XiV3L2JJQKCHiTTHnVom1EoJP+QbNJCh0ajk4lOrhUOSo1lZ57L2YC1016vpQDEaYZMeyHYkVqgK
JsubbCy5o+iIEGQBQbc21DhPfdqxq1O9gMTqyFqjhQZ8X53WaPhcmIxP41/vID87VJ6qAVR59VoD
Chnwyf5/xMz1Mg3jdv/LbuV16YVhRUjkIiYr5yt2Z2DT0lfU4yPmHU+emheIpIpLA+gNRh8A4s5m
gsC2Q1s7eseeVcvJAeofMBPDkxts4p7bR4k3PZOJmRwehaXWYJ3RnUzAm2pJkhvdvYcnqv28xIjs
wBamLa1ecdjCdOl1P6feEDPxA3FuMm28hlHESaHhUdjCzvl2/06yBtlKYG4cBP+Zwbchi87kO+A/
5D5K3GjfW7twFQFZT4w1i2cP4AuMxjtovR+SHevtIJCxFWuyIesI2vgU5bkW7YfMaXFmETVArBcU
XvHTytcKvU/ODqrB4KleOj5RfrWxgWqHk2qLg9u302LyLgof5IiZGgxfWczQZoB62GOujnWQpkzm
yAlzm9jPZkoCBuJRG4pP1DEx590Hm7eiwyWv2a6VLM+eK20uq7fygJAUI5TNK51ZXC3Dh33pr1d+
H4/tiKI3YhvpYPx2tQ10tBb684wOg27nvEFjVALUZF3bEvHn9LjpvPDSJ86wNuhvKafZNzTxOFax
OVYDyHawz6i7AxVdEeXc2Pc3AiO7aFkUOatJQWQ85gaE1/VMk/4wo01Z4PLB1tW2u2VG4XIJ+7/t
Z4FlOLh8iOvgCPm0Q7vCtTMsSSzF8leDtw2fps41a55JnYWSwz5bYe8DFpI5/yUKzXXVPvW1Vrx0
rpoIMjMtXWUEvC5YDHeERpF//woyCSYnl9Z77lAWvawDLaGVWTKflLt5czO4JTlrLbkcAv6o4ZMD
FlA9vxWppEwmGtFStC2ayicom4qB8CRM40V9JhBSDNlOKPvMOB3oW75JbrP6TWyTU8fsltvgXuGo
c75RQ4g2gXz7cigpJpEP+o9aczzI395tYzReqpUmNVH45a1h51QzbQ445sHrjrXXKAKWoEHamasN
4G6f0xb7Ut2HnkwmbLP7y5Am6z1CmQHixvbe76rT6A8bwhCXYF6jZ1yokv9HXDlFQ9sO2bU/x7LV
O+zj6vI3K2juR3ds1jHMdSNnliVPC9guaixMQjusaxZUcH5oYRpLdfOGPPTIy5R5fRkNP5/I8S5h
zw1BmtVzkytRyn3Yp7roDv1zFjJQ+SpjlaEpFNDEMNNYSXbxAQib6LclCi36o4F3b48xdRGE1Rz8
ZCqW9Pktdad8c7f9A93UCexUSBJAiN+xpZpPcqwXB4jamV5L16WtG90f8PkDa2DmowMZPsmhX/0T
UdcopPcvc7+vzNrszHDQd0gtraEryH5lro6SQkiDpD9V6VcnOqQ9dFlkkJEFv/JO6rYU+JTdwkpv
BhO1lXMsBvbsdJ4k7capWfRUfQR1DbpIIez92hnN62JCjpLhWiGt2Hc2LlrT/B2RSI3T6iGlTLfY
bLP9oDcEtkVa3NDxXvfq09z/5dq+jmajwwnZ556fc8OD/XTdFGjxXMFWX7xrrBIwTmXlbFA1gCOT
Mr7XJZ9DhfhjyZrZ1tMaEjreTCYBdxQ2QlvzG+oDUtIRu4phT1Gzg3beuSWnLB91GfUahugqvv9g
CJrY5Lt07/qCnLuVYZK9dLtHnT8Vsp8+5xI0r1SobLCi+xTm9eSjZzuwUhipq+AKQxQEwkXRK63m
UE0CXsvRHrNmQ8nqFkqbXsyRNqH4RS8DxIEGGDLY9cokn+e7SrlXFwi8zqDplwnqt7ALlMAp3NHJ
04r3wRbckjyJcHyua/Cof0ZaVyfq5kyjQicgILbP5M6+tKHtmRk+kXmkbjo/Idu+dF5+4IpbrDle
YtdIotgfYyEPjrBY5WYZYja5nzv6uGdGn+AalyOwsPG0fvaHMrVDVlIPAGhKWFMLhLWRl4m2ww2j
71sZl4xMe7sb12BdxYGCW71H4dGSITRNWP7UPNZ+XpfRYnzuGza7HkeoiExa4EMlH1kwAouTu5rX
M4gj9iCNwQ89egL9lrlu12lWcbOKCc4b0lxf9140IPKGCQuwIfpACMU4PeBbekU35sJnEbeBS3+/
VsIz4PY0syAidN0YVfueSan1ICxeN0P28mqmMUwrN2GcVr4mgKXWExJKUizc8qOtpvnVNZZsOP6j
d+QtjmZWfGkPncQ1WZyNwK6GMKN7gswDGdv/dKFHFqo/Ycb393Gyup4Qqd8YQVqGIkQIIGcuSm+1
6Gn9aBbLP/p367ifmWJt0oKG0/jfJYWF+E45lBkksmctKJKAlmZY0b4Zp/Aa4V2ZqtZ/sun5cGA5
BgMlgk876IgG93CsW0ImcXVi7pcD6Epug19nSBBUVr7/cn7W1lWUSMjx/Qnz/AQhQWGZEO6VGaXx
SZp0C1C8rB+1eYaXKSbJKPeicmv/JVhqcqJ5e8cwi19jQ5rKy/9F4O5pbt0qafFg+cnd5Ly8+H/c
Q6Qrb1NSJ2i67lbls1maz3ZhEbkp5gm/UqMTaVrKeoa+aNJKVdSVZrZhWgIcuPW6Iaeh+7Zx348+
m3Pjrm/OKzr8KdUfKiJhoXHkWqV2j7wHFJu4v5X5gZoOgnhU1JltXOu++2Bk080aIAa7iFAV5nrN
9Sed3a+lCeZFSPukJVzqk8rt6yrF7NmkcOwJeIupqvKSDbcd0tgN5OevWASZTGJaUFUPUVz6UIc0
WlHGL+I0zUSoJWErIRxogs436OYln3+Mt9ULcOFQWAa+ZXWbDwSyuEA/1K8on2zt3y0EQALlv+6H
B2zfkrXg/tzMQUShtrCnXmduXrbM/edU/weFg6rAn+lv01IigkSriy1cOIw0o2SViuBgIG+FeW9n
KIvb0eWZb4zZUSgXZpr2QOerkWSuzfEv41mfiATBFui41jS6LoBxH1MhqJjs7tUMjsCeK3+f6VcO
0EZgo9txCeDIkehAMI4cVRxqHTO6HEbuZMPCatbFxidOqeUoxWt5BdZCic/328IYJp+iSc3vaiNm
BuRLiyzmIWY2XM09l47yUYPWD/dEWBbegw8X47zZv9Dmw2aUmeGmTQ52sQBNxbXyr7nl9UIfSGrs
OHISLNvRpAAFRPaitUC5WZUDawdeFxkP42CSQQazxqt5ZcFHZzo4CUEFzWwOpq6mXQTh2Eek7uoS
A3hoOF7fZ/ILcd/yI2uT+YuI1R+X4vpEWWHq4BaiV7UF3QCOck23gEz1hu/w0HDW6Iebms5IQLvb
oFQEws37hTz0m5WwFjpKc88ybcE9aqNM4CkBTQDgaomOy6H1CakjLWFHgom2DV4wIkzA6TLpnT2P
uTEsmoKcEf6NyS0mIoTP5ZLmC7VcGku3gHyBEWmqL4fOI0s+QMzgq+SzsV3yS46dnda379xh6jqM
3VqvQBzr+H1g69zEHrd2rRVRnwuPSBvP3z8xCWja7STEuk7mAV4pvge6+htuMmYptxTS3mP1Lznx
TwSbcY2B8PohPbqd2XK1fY0M/CFwpK4E16n8ObgrpOre293Vzl7FabEbdmsOiKkyTxjF1DjMPb4S
7t387FRZkvu9RpiMN104h1Y3HW6k5kqCNAuhHbQSDPRAgFQz0sdQKXcCUSKyimBsE1KuxKaMqGvG
6UDX/7GDWs6ruvQRa2jr8Rv4H8aveczyOUjMJsxqtpuS7Q6+uLuM/CrlyV9ijXoWiE3zN2j0bPod
xSczr8dq8/lFktbzbpyQKXRA0XabGnczF8Hq5Geodc0fopCDz3MZn5L7Szx/aE4Lb23wb1aNia/S
uWGFVeDtFesCbYBmjPb34ZmkkeUyhFlzE7JZyHaqqcql4fILemTNSJWDWVUQbK+owFzwWXTfXKKV
DsxJtSIuI8uAgWI2h3uOzibnRzI9qrX9HUL6uuxof/0I4PHy8hA5bRycb78sYlIKbrF/OLHLzPux
uFEpxgs4gkFrDDgUrX0oZny03WdahkCcH7z2NshcIepJVFWfoismns75lN1yNzlV44SVslhLlxdv
Pds9V1cUKAgZfmCfH73KqYNP65rnK6e4OMdJoq2poS4WX2KLTbyCgyt1hBfpczuaimDgpPoYiSHv
5HbCA7NRhKMe2RgadRt81n/ti5mOseH2PokfbDKdIx8CJ3+bcmexh7WqsFYK5mO6r5BpkP4HhCBV
bUroPCaBBbnpw+m2rNc9P2aduLJUEdJ9GIaRW7PYWh6xSRVVWt3hJFRbraMXVWdf0wI8GUqDuVnA
m0TvJUT0QvPJ64YXmGenOrt3hXkBKga+apdq4xZNpu9DWSSH0/jbA1tEQJ0ROF0oY4yZw0EWKuaY
Y5OT8XeUP7E2ZYgOs50EVjXzCN34NS/hBR9rXGvyGIRnvbk9qdKXXtJSxY+w+yV0s6ck5OwY4HHR
NtQmOYALcBygD/IPAZAfcL0SqJsH75ncBQ9GaOuCDbk2xl6b10qReusOHJ91lxsT1x/FpoGuPgIx
CV/PplFABBiuXAAN1aeYjmkNm2lwmzJu/048r07jArantQOHe3Yme1k+HJOlDMqLaCu7L4Oowgly
GFYxu5gqJIp2ckzS26GLPJYr8SJGluN4+2Qs8wyhpj1CNYmC6KJgSP5AesGInuM0DP5FAgVs7Kfr
2F20DgeCzfIDXgfDB93Th1bDF2do2AT/57KU0jpbm7P8Box3ISWc4+/RXHGSmI2BsQF8K9NIhwuM
xkdYGygXaCaqJTjR+YxuCkelXxRu6Fx+O8Xb0bm8ymMApAnbEMz06C7Jt0AI10nRjGdg7SyTG4Fq
8nmQ2Fry6raYZR64DMRtPD77vkMJO4N7Eqh26B9WNJlWAcWev77EFTpIpDuYHEOc+xroapvTscPq
S0En4aDPvfa6ArTESTv0qxT6MeWOu6tW7iZIWqUEYjmHZJTilPjyiEdFDQmAop33jj1PC7JEHdmS
9Kg5yW0p+xYWSX+MMRBbpFtzg7w1J0+A2YUDY9c4pZ+p6v6MrOLXoLTiIURpLXM0adqOoyjh7HuP
rKzoqqsMM8DK8ClH6uqsSC5iPRCbGnO0AgSAN7D4WY2DWff0gWgB3qsJUCiE9f+TxZwbaBaBfv82
dLrCkNmN70JETSyYHHWp3x3CE2VEJAvj9YaVQMyT2OAFr69m8twNIuQGqIlhYgUZCq9GP7QKtxS2
9avgoyMhKG77ygOW/CP90DBfVQTfmWrcFGeuvEyAMg399NwCIYc+18RKcX7TEIgzCL2eO4lrEJ6+
FAUoPx6FqMWje42WWQHSoaOwweYERWftvImb4qtBIgUj/BaA5IM7VshLv4WbWoSgcIldai7oUAB1
RIxtSoCwv5Vg2kCqt8X2bewwPUWyd7fN3xY2xoQ5YwsHygs7gmTVnXwIQPqwtQ8s4zVYknCji0cW
8/Q9fy5M7lIHTpc6XBcwxpgEyuPjDaZWDJ8mAUFf1eHuuGfPPjb9B3cyHE13dFvofw+fR4EXwnQ/
ktF8Gr/eG8cD7oXLSOgsEwkn6jXzQluX1GNnRS06w+IrinVa/0taVBsehJh+5TFMKTdl7EHtUv+n
W7ECR2u7Qd1kgiIzhHwsvHW4oWHYVpgqDHFOEZUyucgUpt/kjLQ0tKwPX73xWsgof3wwIC3AdIxh
RUqefkuvSDCN5lC38mPqgNtWNIIGd5a1iFOPKb552N9Yg6VhjSGOesBZ3vhsMs/V5ocIsRk0bFdV
YsfASWvQjGGPRQCQc4vVHXirtSiY4+C1pfN22UtKVLeW+r0oCiNV4n8lvsrl1XmrZNZV5V9gofam
aFQqJt98mfMLr9ETnXd8LTYq/lhnBAJ0kf40kNx8hmAjNoQ9jZyIHJuS2lOeDGI8FWqHvmUHEBaj
Tw7QsiNQNjmGNIS3gAp5SmFVu6+KKO5kiDThhMSdRwV66uMZGF+ZoKgzrKuJKG2AoVllclT9dXDB
sx4apg/AcD0GDfk5rt9ka5W2gyMXMdBqak7W6hHK8mdmHJ3DUETwqXFAGqPe92AOS2INW/ZSO5Qi
gatDdo1smc1tbhuR6NgtsAC52fTvUqFjDB4PvFdE++bR1WEVAu6OJN/V5la8WJQLoTcBqvP5+Ucp
IpHiXTCsgN1sevCnomkVtYxVxdIm+aca596nZZXDFJlN7P7Vq0YqRfhUQEYjudXb0/b6rzKJZI8B
FuM2EGXhDJnNnW5Rdx9cFk5UaBIB6pxUIVwQYtWQvpfEIhKB5gHVcjC7lVVCVtc2pPsbh0B9iv3A
j177/ugxdbkfeAtsM9Ef9Uc8EjCYLDmMK5MAKNGSRIMNTv6/Kvj+iDL2IiBUWGUZgZz67tknr0y4
Xh38Y0+qDIX+XPiSVjwfXaT9KamsH7VRsMMw1nSFax5l8TqOkcT7IAtZxD2PRpdVzGIb3ny7B/vd
8NrnOylDH7Up0neQDBVreg5Z70GK/3YeEdhgaBv1uum0+RM8Uk/er4cUEBs8xtNzXIyiVGZlciBz
gpU+jj+a/cL1Ju17Ca8UNKQzBwirtC36egRhTrxG8LuxxUEkBM2BAXrbf276AB63jEBhm/mZ9T6/
zfo6FIP/Aw5yM+m1xT8pBWYULxkmaSJARZIb0zAhv096Dc5u9jkhbkjuj+xZ4DDM2zkBOcYBc+8F
nJE9T90kvFLDlN5ZOsRGT2YfXH5bbSZsfKRkXPUVTJpxfZVVTYPXNIdbOT7rG+/uqXM8kt+QFBtJ
Zooj3ZGxUObxNnj1vZOhQGO6mne0RyMeiS2ARWRIFEttgtCI+lpBge1Xs3cwBfNrbnZyizbD/biT
wDzwpNg1kgK5Sjb23K4Vtp1g3r4cGIaTJrbDrQqbdJhWHcGYaEcN2/i0pvoAtMSxkmQc4uFa4Eyq
UeP/jyVlJE+mKjx0a+VOPc4nLm/Av83XQui0JR0tmAUB3bXS4hovf4PmjS3Wk/P0JWPUmpQJguom
qKYBwiGBS5azDOSi2035Zyw33flAs4s1o8ikvXAUTtG6SFWjWcQu99PgFs4ux4P/ZGVhS2VriRvO
Irf3SICAbu3j1YnrtprpL4qpDpYZ8YxXLn2klqKQ/CjpNSjhhGlt5ISF7HAZkzdFh/mlFNYMJFD3
TBwftH/BLbxwXdRHs+3gn8bfho9fC36UCq8wYtwUFFJDcJyftyRDeAbi6GuYit2eu+kD272wqGmH
ykyaHnKRTRC+iEYknyRGCsOBsvM8BOPMYUe9TlwbneGUA+cYXKwq7yltwVjHGoALUgEOECjCfbv8
pbL/uDI9S0OjFZKuAis4k03cIf09PCpL0dhONBvOhpJCkHAX36UWo5Aa1ggtizOITDeEcKn7S1iE
JsvRYEhzud2qIBeMFYNKcLgN1FAJdzvrWnsWLu1ldHxxK9Adj32u0YogSJNdEw6YM0ef6i5UZSjv
bIBtNqMY+xcxSGkVjhTn5fRkqcqBdhdMNl8XndbXKIdBH6IhDa5efDSk8XH2FM0WhGuPjs2AyoiI
DiVV31kH6qjJfRK09XiNXvS2DYkwAqyMNbjRtdEWTle5Bqq0XWcpZ7KgAHyKp99owlqaKcYIVXRE
jBHLQa8O+H8dwXYkSCbimcIatyuCzFIvPiCUTOITXEM62nySHlSr/UU4mMssSBpnMt6hLYg5v+fD
ny5z4WzzAOgPjKIcOXRQDNtk1+airNQxPPLLACMZck+QmEe7LCTunrwUauDggeUcx0cdFwEFAF32
30VFmggk3ZoTxoquBVKhc56NrL/IjXFNJ0Pi4r1sgHHDq4nsy/4fnqOfAyFv283w6z04Q//iuX7b
thIkPwEhGYs9muMyiqapNzFdpnPPg2EzHED6+p17UiYw8iJbHKNnfu4pAIne87KUtkl0vyOsBxnq
wRfEud5SgAcPXUT6OA2lI5jlzpgAozBS+3Pkd/4TkIhGdyTKaqso2FGRPr1mP7Q5tUwhg6Xh+8TM
LcHxSum0SYdvTIYOeGZwZ+w0HdDKKhYei1gOpYEaPYjD5E/wferEwkeTD1P8CBVVJaiFBk3e2xb1
XC+9IdFo5wls63NBocxHxd0GRByzsQQHeUTg2HgpuPUVfWV9RE2Vap0xj7iXgX/OAeJ8V7a++YIA
ZhImjdGiEL0zuomL+Q1g4o7HkWVJ98MNonR/ITOh9oP6CibPYZ9eiz25NhcTvct8q/4gFfLGSyga
m60OsvJl/orFh812Ci1yyO06S7/k74cBY2uaKqit7n3k6wb+DGmWAC96Jb2uG0gEzyZJam5YB/Mh
MqidCXMMF+qaE7WwqbxdtjipQdc33RIyom6YF9OmC18TzPQZuy9BjgrghshgLlIuUvf6Bya0RQM9
vqSkV5CJrkobhDheIPIR6ZQZN5F3TFICXT9KJujG3GuO8KlRDFjtiW57wjjF3FuMnk6qqzWho++k
C040WZFh9jy+RuRrWy7bHrplGpQg8Vly3ycx9VYnJDTyhnT4zzuk6WKE7CtBmLCBRhz/y/QJsDMU
QXXMlle3yKLHqihZghXmmk3HZ9q04VBtCmVj+jQidyZjwKhcasF54n2A0YjlTbPxxOlnXI0Xzlu5
LkQYoaG9jts8efrk2JB7znunLip21/Xic4qr4EgLB9SIYfY/L7srvi/cPloIQrRf+aMKFvwrnd10
oDGJdA/Z5cfuiaqwKiZcdHFhRBNCrKZI8SvX7DPVtyckLep8d8pYf4KPA2uQrbMwRQowLeq9IihG
Z2wgaY7qBgqPK5mRtGaJYnlTSzNxxHh1sqI9Uy3xgYXZ2Tv6pvs5dsqdkQpiD0TTf25YaS55hmgT
219cCZeQ50uaxWPf0ejYM9wZj+k8Ktizo4p1qkILwdiVT5wphaxWeEc8PAAUF1t6jnBr5rXPmBBN
GoKsOspqJyooLVbMBG0t3dOcjOujwqirRnmvKvyFlMuQNO/lpkvL6s+YWyv6Yxiqf4QO8akkUy1h
M4tIEmMBkOXwFtJXen5mvMRWYle7hq7GA1fBonKFlOglNVxBvcO01pOJeB21vOCzkuZd/miRjiaE
49kjQmVncPt/q98NuQHeu1ccdoIOMhIxQMoNmvxRfCAqKzYJuIGLXVB7QJlbjX2/N/T6c9SU9+Cl
2l/3ijNYhTqbQmMFoYqG5fALQchXAUP8esJgmFZSbVdcA0F/jzePtqoKfqOZifTSp2sONczFausl
5SVHYTBsq2rK/byx9Dbz5/OhTOmIeqWjdGi6TtLTMO/9SD724DU4JrEe7KPOcVy84wPi/xGHFROR
lC60da7xhGLTjMeaCQHwGoJhVssMD+Nsk28olUz74+t5rtIAH20aEEklsSMdaIYOargFRgjLjGnq
lNXM/2p1KixJ3jG/W2yStbcmTaKnXN1TLWH2/Hz/ocGMbuMhKHFcB8DTRJA60OV+IonVljCclMhF
nRnoxWWsJfhjrPgKsz1MWidCDP0+jMyNyLTvdS5vGFTJOzL7TocmjG0MdQeNErvyo0eTnd37JfGo
Bwhiz75NUq2ARn7dO1zT+0/xLABLXK4WXTH0W8g4qOvcG1f0tPevaUcq6THZT9pGQwNIaBp1d5zx
JcgDbQ5zocW2+bjyrY1JFbiNU1E3SUXXsKgVEoUxQO4lEiBVBnqoSjErHtRYVSVxwHK4q6fqPPSz
SC2hcd4UKq7wJT7nEEe27moYkA0tC1rkkIhtFQza4t8KA8YcBWkGM8uEjIACzEfVjZPGxZ6B4bDT
e4bf/oUUmGvhWsB0Bn2GGtVO/DWF/pdYLHZSi4erRvt2QeoSNK+8Z+1POuTs8D9dRUkHqSHnpagT
56rCQWlV94riByAb2fDmfTzXTqFdk4No6jV2Rg0BnfRtrDKGfstwSVGDS2rgnS2uHq1/aN+st3fc
ONhfYUXKmzn8YcSLxU/g1dfNdnGrqJ0JixIOn5GmqQhlK39jvI9BKgielYk0BkHjRLSfP31EgHTJ
MAoaBxuGShki0CMNqzIXZ9xZGp3P6bTl9jtdxYVnQpyghviRuGpakwajyoJtfteLcqszZdpH0/nR
HadkIKoghiruyq+zuQ49JtEcuN0tWYKEQN0LxcEyAix/r7YRg03/TfWhm3219/jz7TaLqV/2gpfL
o8txQPCFmn93V1rquqD3nunMMgVeZ7RRLGrVGIf6xSoZMsTnVdqnb3OMia+5lx61zjXRPbzyTbZo
YTJl87NaIfiRA+yEBIFE9cJaHdhl1WzPGCKHLt+yZuBb7lhijyq5CXL4vOtnLK21AOK2Yhm87WOB
lw97ZKuE7x3LU2F/HLVedl32P2B31qPtgDuM8HVdfbjP64Ir6NK1ScVl2m6bUkr86sGLnJwkhhED
J/JkGzC8WTakjFQ55iBIWNyKk8IyOG5ituxk3N7Ks+koMY1sM4fZxq8zW52O7rCWDXAiQDbAv/1c
jw2sUWzIgxrL1lLbrB0J9yxLqDEaO35NkrM88eW6nuBYIxpPmruHo92g7fGwGqFqCAGQbqBO/245
QuWAf7dbKhIMUUUKn2GUfEqIZLzkEXFACZHO0mEiAPv8gtj/DY2d61FYklDMNzTT+NM+tHOan/N8
fFAj3AgloakyDH9haGOEivYRQUIR0R9RJlad2Yap9PrL+5fxOXimFODAdxC/9dcSE83YSaRbi4gs
uVcPSz1G885rts84WDXcyrNStcFcLovPwGz385lqvQEvLFLEvH93PJ3pzZOSWnX/l8YIDGgSuvBR
WYvZ7G5o2Fi5KHA7JBG0g7mgE2di019xJn9EAAW0EFDnZ5Er3AZi4R9aCRYOoLX+spz5AeCxRhQm
6pT/9zEBur1UGl6MblzIY3rDJeCc8dmwM2pTIW/cJlIQBSOkV7sZX14zeDq7cep0FQrynpQxj4aM
SW2iSqZYv7Ilue1fdE21aviV1AWEWLJ8nbzAKNY32+pY2YUq1Dqi4y3LD8/nEDnSzMDKi2t+yv5W
TqUqnWFRnBxxCShiaMozQ3VbrYF0FfcUEW+qKbD0BtltDXBGIkUEEEwyD2TOTokMDJHJyltq1U0V
jWmhvsrI371Pq+7NyIjKsHApsMBveX9IUGTpRa6AFppAuCwnKdtU9XFpmntnItHWAOH3QGBcRUBs
4SIXLaAUSL3YJ4QwoHjuByaI06of3n64FjRKO9aB2Z0ozdpXyXar8MZgD9CbNE7I/rm5EnHkfRux
9QsxcrF2vkx+0qTgfwUZrqCuU2HBb+MX8KKUYQni0gd5ZGFw+gIEOx+R87dmZEAx/qTkfE1AEN0x
ZlVYY0APnDXqCSVVx0QB5Gs5HfoX7TW8Au9R9j+bVmRl+u82vqJl8tkx+bPJzUQvm1XebsrT5fjx
t0t0NwpYGw5F5UHVzVkvg8aOol/L5AuG+UZOk7wmTRBgDIEX6g7B1yIAM6Li06++QdMfBErZ2O+x
RKJvU1r+xrYQRJdol4iQ2t8fYJeyHM2QKGVKDwz1ifMGKAthm34lXSBOIcrnQ41v0t4AVPyfMrC9
iNan/sWbHoWeKkEXyo8zYRfk1SzW7TjfrzJe3gwJKe0wfEoxmv7c6PiFXgTVujIYwmrSJRHbPMnt
KY8i0NkXtMmd+KYJSl5FlyDtkuOTakLR5Oc42SK0b6qAnXxqm3PrxqmOqvhEX6PlLMGhrLQ4XgmX
r1NvgQHzt1n9QPJtMhkJSznpAf0ipEnIECCwL3yEkp+pz4knYVHoXD0ta+8fQeW57x6Cb3EQFE5z
HK807wUSR90dq+fuozHN9Aye4lLMlFApwbjg2r3WstFn6c5QQK3Yx6KHmC0vFGSAC4zesmHpAU1C
mzaiPCj6Oy5CSbm3rzjPiO6J9+12bjAoBCI3REGgRgqnpJ0sQosGMP9EJMV/APWAEK11kFqMcHCy
/vaed6yKF8NS1VrUZFBDvgbIuLnkzek+/t0eicZOwmEM7bRDjKDvQcUorOrPoNrSVvgSLAA4Uh5d
EjU4+638Pmyf4zcP3wB4QmS4NRu/FT8FGPWQyT/Y2K5TuL8jK3GeI1e8cTMN0yimh6Sii1+HIuOD
s0vprZx98qsttZS9AQDAYvhATT1weBx0wAm4t04l04KxVFfZ6jkKd82fJ7ehBLgRD1nzBsnExw26
rqNlf8JUCTF1qLfa0+JS2yMWG6CTDGQjZL0QJORDjT7OneAEHdKWsqQvmbQYAGlYd1fOXPa5eqv4
+JG0zBq05mzLbb1aHp9Uqci9W+uDGVu52TgfcSyZ2On5P5WcrEPDOK9gZ8A493WWRZoR2F7Yj6q1
Z14Iv1HzKDb06S1GOWpMIgg64/d8O7O03B0EsX0RphoYrXlMb1/S3gI5oK66ipy/bdu5q0pBABcD
/WMzkMnyTbqM3waaMBGM9g1GycIe5lQamKZ8cdcqVMLZzjSJTi9kgQfYRMHRJ8LCsAO8HHIFpIER
XZeJG+qYzvCDEJe8xuLlj+mcNElF1hRhIbk28Qi3ngDkk0sMSPFxpHn3Crn95Iz3PTFv+/KUgMYr
WSP5776CAfCAagfw3f/BYcvAMxzDCXHKBxuM0o49SoRonEc6ElaIZIo6/rokiLjrqtnHytU1ZGj/
pTAnj9gKy6/7ep0nenxqc/vUsx4mhThciSEPiSk1sUOSZF1g3Rtb+xJTDNQoRMcAu2LLpMtmGkVl
DMyAVHOXFAjuLiUHAA50nioipUjP0SrU5G1YEQ1fcGTya+TB5IxH5oOy2V5bLJY/JEbByNoLkZLH
Gafn5w69qgeK7T7U5Zb7RMJo4mffjK2yP9gkYnfBZsTjR31Vi9YdkD8LR1WBl5mKGLTbDlyKiSLk
LLS+kg+2G0d8iHdXUAc2aiCJLG8dnemt+XZzCitVBShFLRfJlM/fWoUX+dqFCg+a6OgRUxW9L3So
A/b/ih19ZPKMeoCTP6Zbd4/0rFzFlLB2mJNZYXDb/pR+dU3uRN+MW1gbrz1yXlDmsVTQwaQVvsmb
5cnOaV4BnMY9Nx1f3HWa2Q3q5tVorm/gBsQ5LixqXnibtL8xJdzBwzUCQN2CMq1nxTtxNAcZtPW+
au9WBQl1qUdYEPvT29K/y0Su36PwHbRTqohOwmJOVsaFFYraefJ/59bAymLxDWcNIwOVVfi9HaTW
zbuMDZvGyyG6isCIfXoeVYaAd1/ioQI7/zX7eUxFvmvFdO7DdIxpVX0LM7q0IR+/fKcM6AcvZJh3
xxx9H7H03H9NeLVocHKZEzBUtqen1uN3iE6pSqpQQ9a0Vh3G0+8DgXoICPS6tRJoOU8EZgFgUd8i
dIqHAHVjUfNgiT7dyXGhasfP6mCQ3PDXvIWOKg+a/7PtgSU24PuH7p1bkNtzJrhDhLJp/mAw+0Mb
HbKZPRg/czgQPPKzO43fqJykoMCpSCNwdHBGGQgRPYfjjx5kyG+VaRsBTgqU0HjpTgniSPbEm+94
Q6nwpryaczLemwHKvHKN2tZVri9gsXDTTdIsGUpMLErkkc6sQRD3b0pxFvPZpjfzdJU8cNao9F2n
iWy/qbCmc+yodCkyhXqslF9cmh/EzNWGJP2WBjcNkNSsUZhyJ+wo9uhsn2wsp1akyu8+oCrqoDkl
7Hea6bzKcpoYE9IUFpzBxI9Qzu70KEggroRVqfVSHw3YZ2QsxhocMVsWRBBc5XNHhe6e+gqWZR5D
wQ5lk80nye+Ap5SaRwTzX+Eh3d54GUAVxTuEo9UPGahTHunQEAhCHoAow4KJ3JCXtoJaL9vKja7n
OFuj9x8C8mrkjwIvAX5FCnsNF9SZ0NKodlYg4YgaPfmmUbuyZ+pwPTGgXZMCQXEPZjzX0cK8oLfE
ox9FfsLBCDEhV0ebmMYtJzN9X+el0ZwB5M8znY+BDoArWDw7NCN6FvpP7zXeiyRMh1r6Ip+N2SOY
x+w3/Blx2B/ilq3Mcr52TU4TdOqRt3Ovu5XxE/s8xReoDAinh4tF9rhqluOuWpMu2s/zbJdRQU7h
TPZ9JqvCVOEIZ4NbapS0h/kyko8Mo/NUN9+t1sR1DA+3HXOv6D1T4W3IGnkIjnx3gYvfu9bnMl4n
R52H+thy+gDKfIbdhciLTXzUtvvM5ZxVno2usrFO7wD/Y1o8yAe69+QtIb6I6gv58aLNW3g0A24c
56QkbORA7Z8e3yUipn56PP3iT4ezVdxsK3x5RmNDkjJufe9PPUq6DinzQZqeMOf60NujTIFFSFCC
QSZ7OJ5n/socV3rQUNJ0UT4W69CO2x2NpGqKEGACp9bFMTJt+RddMPtbD3cxUFeOA7oB8dFJcnQn
giVbE46H7ZzKJsMRp0Gu3iXZY8vQF4AIuK8RM/2glj6/+VGMSq3+ZEVq5cnYVm6cKF3qv7JnIHPG
JldvuO4cD5shUeg/RiSvtUe/TeUkXuFl6oiSFBrpZZ5GDlpQD0WQ5HTaNMWYA26EFM+b+aCP+KqZ
guWq8nJ7eVPqfJPc+7FxLoymtlR/H3/qZLdJW7Jfe5+EsoS+yDpYtro6+A7qMezDt+EQkh67CoTh
2726awy6ZhFGyH4qixBUZZ5gKg9lJZfX59hacS7ckvQW2jchjtiUpBOvk/grfLO/reA0K7EjJqTE
44QxqZq+7KjeHFha6WUpGZgQgkCqQi081HKffQ8HAuCHuAbx3f26NvodTfEBEfj9jSiPI4ymRMsF
ERXeKtcc7YNxBK4BF+Grw1Zl71MU3JwJbTNCSwMlppZyWlklH/odsVaMiaJl21ijg6CgajFemN/B
F65v9LdvrY4jComDKIOBiDrLc9Z3jmnQGRqm0JIJ6voXrha+5MtBknixmV5gLFPzbCBkM92UsLnE
z2iHBf4Y90WNtwrX2QUrfzaoh5HSyw3z0YfMZMp5DAUJY5lvLg6ylVr5i5Pgrz19LwXt5cZXxrRN
KhtYZpGjWhxiX6JTpIxXUeCeODjT9KOnCOIIBijWgSWGjKHrljvfAb09evDvp6IMmh4xUFr4Lx+i
4oBg/y+k5wOKH/KcmmJ4+nK52MonJUhQp9brs9+AvhDXd/PunT5esiHe/nwUF7VD8dGKfX4ffagz
pOMdA+oBUwIQQ5yUwQSQEiARh1rTIJKk8/9JHi+DqV3YltRiHDPs7qTSZBJVzghSxGry7OSjgDtZ
YMuXJkWWeB8iezYIMlJq717q53hY8UvOYpJCFYtXwYdACjMwQLufWzp52jUovQx5H+De+0f1I8tB
FtuCLo2HZa7o1PhoKUTZPXLwxfODbJG4uoAhYv3yy/kcnCHA9+jivaJlW35OAEZKVk7+Xut1b4rT
1avjUlbFx6BkVjiI3JLe7nnqRvELJ8s5CljRJpfWR981rJ/QnqLHEabjOf4lbrHYTzu2J0I4Z1iG
LDYNvXTnZnkRYvETtmcBgZO9SScVea4ce944NLbX+YV2bos6Sy4ClqLjkd8O9l2Bgk7NLqidk4Is
2i8i4bqAzHLrOBXU0u1+mu5UmLW1JJaBIy/D4znjG0fYzRE2VnaJVMhHyz4M6XrGedEp7te8XjFm
HhXpQfP+WTpH6E+Ksv9bGS4RlSXudldyPkK0mR40nkmoFkw8jTzhV2mLvseGkrVqT4HZ9FuN9Lxk
Tn5XsILifI9JYaVRRdwquBYnE6xFdz4X8ZMR+aJPPtrS7uWRg4r5PouPhrLwIelhZKpK64bB/o8Z
4CKBDDm3xVwENv+MqRcI7ar1+ie++rHqgQlrhtP3AFRUc1/1azYVnpf81A2MY+ITneHvaugUhsiH
YuD8q7ksW1QCTw/J9yDT3pEXLbNEDhSHQCC+qIcIQEwBdaFuHQgc4oKMbuuO17lear16/7oPLgvE
bcAD2B0uSTPL2oe1Wp/+Qy/BJMomjb5PQB3ORFFDEZ1dkTynFZyjBq1zkWFfkTGujlQ/2S28q9q/
6EEUkC/byrKCSLTO1YZ7hpIDcSJN2+copk0VVJJ3MUJpGCA6XS1b1lkdxXeN+IaEI0zL/jqk4NWX
pt1iSzCKg+Slx+K1xUi4WK+uW2Qxcz942VBm95GZp3dPOF8NLr4aQ7EKi9Sq6f4/U/wtpdHXAvOm
088sBqCg9jDWPEPUVa9AIbHJ+78+RWv/z4tROJLUSqjiJXVkNxJ/eV76ngE7yrCTdeaBxNANI7Dg
E7A166l8+5yOXsHe+CxcEFs+c0qdH/Rt4K7NvL4bJx3bB3LqDke+KPP1XBYsxkVh90nCavglAvHR
FWVKPOfaWEJr1q0w+9eisIXyClwWgaIAZAROtaFY5U+XKH9xm9YARvAJ1+jvnRQJZ08PNEaoRqiW
meARUxDvJoJuZnmHdzWX3wCL28ybLaCDRhy1+Z83u3be7zzDhO037jMHuxV982otXqUaGwUzvWUa
3S9woFzUOoFYIlQUzZACv4I18fEsBvR4iv67z4J7nBcN5Rg3x6oSnIyJdNgh/GFZ5hDKokMfbvt9
dAC/vC9PqaJMJXz0okdn6ktLze73dpL009GWAl8ZQLHVCSxdrjTGUe+6KiW+DWx5nK1BKooiQi8W
CO+1gTLOpLA1QRdm/7/6J4EYFCCrEWRwCi3HmUFdXzQ8xZ22lOwJdHWRmzR5WX3iXwInZv9Ot4Tc
ajOHl0MwMGvQ1Iemk1CPaZUORkZmhlAV7czoeLQd39gFDepz9GygHBGNY0qQsr6LMaj/UpSdiOvl
TqP+vkFjuQcBZt17h9OJEbBoZb8dh+irIODjwRUJcn3XPqYDG+enrutDQCMkIlclrkEFLgtVbgNq
McK44JuP7fMx5hOQ6ohzBuR5nqahLN3JhuMpA5bsCiwYopJKFMi6LSrjlsQiO10WhIWHSyu/cuRu
7BjX64xvsBqRCiY3AUnHP2Bnecb02xyxopRvhnizmEiof37x3p8hhXNXOJFNSHnc+EBhcmdMTvy6
eO9Q5Rtf041u58b97yBPxxMd/phMvb/5HMhlyFW2zmC51Y2nj3Pz5lgYlyZEN5BO5ilzgXLs7V5q
lQWVlnW1xLs7x9l4aEHpsRr28TB/sWE3Ox6tStrB1mBPDcjE7smMl2eHKaYM+jFna7zE3KLSUzT1
UvM94QmNTCo62hTJblIRJDTAJeFEcbttRTdW+o5aYUQ3/SctTABqPBorIdwGSR5FZR0HK8XOu8kA
FjYTt3vwBE/jjed87VEH5rZ96NAvAUuizEoFf5+LeqmCSglviWZim7HS+wbaQbvOvb68plxlbw6r
f0riMTJmhT8w2F1gmlTOSWnGmKP2pQTbLNPYF5mCAwTIWyKipqoGjgoJsRlKEkd+I1F1wHjKTeNW
pVkx/Z5DL4+A4ImjdAJ+kMtovNatIGNsUbpPjdh/YokmX6QRA6qgAlpPAzh6JgkrbDePze7Oztn5
tzimmBwozHq2c5F5dGNDzg8xC9D8jLDq+s3QvI2Og+cxy2Es9aRzdJfUWlzUGMm7BMSmGB5RfJcR
3F8egHmkgLuaD7Oc0e16d35MIq6eumcm1UpNi1i/XuzugaYnRSIiVFWMI/GAesIjtFn0nep8EWNf
dfUIvJGxsM+PNGCaCfpnqPEwbG75XE2nqusYjXn4w6Gl3bgcotr0j1K9/G/H5UgNVaatWef67u31
HARgX6AZszJ1VGAsOaLxPqGKYnHSVZfCgnZUmvzUjfQm+v5IU0gWyjxOekAyyORjH8pW73vh+jaj
ltGTwBBxvRNZzFVNcAnGBVd7qIEfYHjV4ITpxJA6luKiBb7qe0KL0+CBAkp2QIiVFUdFsIz4C+RO
Aj0207GftU8dR0WskPVFUViIZfZQ17mbN2fjCLrDw1TYfuW4YP1yCt4Wdshf2O9MlU6lAJqOsV3n
yGeNHOcfqd+/NEZfPs6jNneaEm0gdAfArMytbQTIwComvrhjPt37uVwJw4swS9Yu4qg+k/tXH7nn
wPUinttvf8/29EGP6x7g7ib3eHUGA7Y6l2J+4D5KT7DILqlFMzviQ2ub6juCPG9+qbJZ+KQgTVu9
4NgHldIeZuLtt9Z035q6l0+IjL2+BtMTARomaV+IW0mdOD6Ik7dP2rV8LGboP6mEbiFYEhO1DbIT
Ms5H1ufClipyeqV/a6Sgq9HVUyUtA13LrtuuvNO87V1oTIakqxSevJcDUcLbTJBjNmE9gq2LIeCv
3SvqMAoXoK2n2h747inkPx/WsFaJLT7IZzuP14QYuE+LKPB52H48BvsXAtT4ER24mw08OqZ05SZs
Me7JDVm1toVgqzDmkLiuUrUxfN0cAr/hZFmENq0KFoFxc0pUYCq1cZxPDFFf74eMcg1FRsQBRDGc
9hck3RbZriWql3vhPHTltEF6gVIUyIHtXgmoPRbzuuO+Mi6gIanP0DG1UNhapVv9ipMbJ/rTIv7g
Wj3p5yvRPTBRF9awMXxpwhWepjTvF/ceBuTG37U6PKf6E7p+d7o5T7CxbMZO23rdm20IW5c+InZ1
FEWQYLcuGwLUlOs0YXXXQnNOEJISp/Bphm3hEVxKdyf5t0Wb+3TFG7Ttf0PAB/swkujDyH3a8KfY
S1XGXM/fne3ODssuMSQZCyiCjKpQ7ANlbYL0NbtNFyfXgGGDRpgaQ4QWY+dx4TP9g0VgIULA5hi6
1DbjRQJCSWFlX9NCNuCjngb0yFmoSt1BEuDtfHDfTIhVqzEKCCxAKUQnw0c2SQ0QxIS7QwcaRiqc
mxO3jUi9US1f6U6ujQWd1eexX0/NHSnOcswDe+nb3RmHGsmud1sJdu2idd/YhohvpC+cbACtniw9
6M+Zm0IbLSL04cmklbt5EgMU6xglRePwuyU9Zbf2sTnxyCVd+mX2tAmbbtympYBNbFQOogr4SP56
m6oiySIHt+QIG4smAntB+dHSVplGxIh82irYiKdcE64Xjbuz6pgwjbWRph182/wEPil2AT8Wanfn
U4gjKv35Q0f1XkMS9M6YtKOtGaIhNV9+omvCg9zATDevYTZ/biJQm4Eb56PNfqxO+9GuNWwq5AUb
X7ThQhQClpPs5jyHDLRZefK58M1t2mN7/wOXMeMMfZAAGgWxHjjJ44KXT042rmGyg9wpab9ZPBlY
kL2istPa7h9XWH5i9w0XmiWAanyg87+N3o1+8RKaY6cI3Co3JeFlgK/wtg4t9jEi6bMGKxTkj0uI
+T1bH+Svy7BACeujDzQOwPYxj/IfnXW17JT9lAqW41u67Hz3SFflsJ/0+bSpa7YP9iIXCC8DNdDl
Vnjh/NK6y+8mBA5vCwlUVWOY8fD92HuKSXJQGXy/KGzx9b/CJbJOalBykv9hj89ZZendz7OgmFNC
b7hUyOApJHB0R+81iF8l9JIcEmP15tTu1VIqNJnGj6iiWxLCMdkKZHNsmk0YYrYcCzODR3/hW5Ga
idD08eXm457vir5QNIsbh60GDcA3E90O5ez8CxJzfvknrwT8BokPptYveIdTJEGhkR6uOzXZbRQx
41mahaPjhSj8u5u7YL0E/58APh5sWPfXbdtmnHlQu2SlGKQnNwn4Yu1uM7Vm4P+fetujuqKs+Qfs
808BXXXShVnqpALGX1VQGA6a7y+c3XTHWc6UEPWRERNHv5YIITaKsPmoB4QteqrzK3hcD6391Y6j
cJTEgc0kN4URtIfL2lHh9vIx1aylsfFi0YKjYyIfO4FDa7P/TQ8bfujRHgnM1PhWAiGjHg6giUmq
TN6+ezZYxz68zy2Eiu8conlLuy1s/rXICLWBAk5GTWU5VzVUr9zYR8pNqPSXBM8xWsytSE6NCe7m
h5xjeEPD6Pwt2mlg/hYZSLwyZSBVyJiwteE1ueUJyeS0fPlFF0kqlTMmXJUnKQqZM5gWC9QBW1nh
tsQbEbJoGM2WnOfce21lPLqyf37uTgoZtUS8Cep06eOz/Q+BGkZ8LyTGtkQeXnyCH/YggfJfNiUU
DXO90GCaTbSx5oHXR73yyKlTjFOt8l0C3REtzlUdWivkcMLD5C8oJ5auWICCHMSolcv593il+hDQ
3bEMjlGtsAvm+o+QA+vwjkEnH3IW8rekiBl+paxma3jlI2yyWHO5njzlk5NxZGJqHZ3yUYOnARki
LgDhb20aGQusTDUizWNlp5URl8w3V9m0YddXRdqFVVTVdyxm48+dbczGB2QoYWpZ7O1jebWgGZko
818jD6mwv7+xMg4LDzJcsuQMFUznbooqHc2DaeW2CKPnOJOU/i3LxqeELoTIXsqNU9HV+k+GqNMR
yBwfrxWfVDkJExiwFUyPSAHmEZfi+vd15fV2dJsQQpy6WAu4WoTj4MMWi5OMKz+MqU7eS9zayaIi
fmx+dYGyDbU7h3Ch2D1yIAyFAmsoXcuIjp6nsuJJ75yOw2xiA1C2lFIoz90bFFcDzubSOzXBIdeF
NFz9MZPb4wv4zcgJjeeFBzvDxgjN2KFnTEkON/5CJN7ea8Fwhda2EUgcQ00AER3eb031n7T8t/ZW
FOVh79iQHZJDEX9C0Bg4bl8fzlhbCIbZlWZpE1Xsj6eBzTy4M1QNTAhc2C8rnC5FQ7SJqBwfmCZF
J8Aw4CHDH77mPqTzxgzwL9NQWPXxcXjmiLydLmrLjvab94WsEkmp2DjpvfWvX7uRsCTloZNJY2O1
cR+YYe38dZMZuH3MAUwsSHAak9PK7dz58m6rxG4GGg9zWWCSRhypQ8qqoQeKa2MQlxqdoNe5wQhj
atWS/NRicvyR+NYp5B5w36WPp2cydx80sVkEttRK3WyC3g9x1pAtSM0svrTCxmAEKSn6kokFDNBe
ji/+llE+CJMHYDp9QDnrLubAcOPPF6/d1Xo6LC+7Vkqcn1ceeBSg09Ii6NFLiGI9qNQgTYTn0C/z
lKCpWleCmprwK6jG3JRPnErHM/+Ol1SjDfAUXZLRBtwobGot70bU38x5gan5b9iMp/epbWB8mH4P
5JUZhG9CWV3HE1+ksWn8TUIAl6Ec7aI7ZBAaqu5jKsqNpBXWBdRd0qmvtJ2I4GFkjvPdjvGsCDPh
6d6yl5NJ075CPd0FvwEmQ0rKJdF1D/ZSeLLKNm9cvF9W6QUavZwoCtPAC4QWFjuOneWvE41CiVKi
3J6YKs9wUh7f7rctzhqJutbMz/k27KSMm+dsLoGhwj5q3i2oKpfeS0SDsKqkszlO+fbHbCal6KE0
K4bgVD46vMT3ASHjgkruzyjY9S9krdVTMBKPhcTEe9Z7LctY5X7+yOVyriMpwnjswYYvIv0FyU2B
CU+vZBSW5hhLmR5GOli4wCDzSKC5CNJRUdFTjLe8oqJS874EEu9ou9/4UK2O2yYvY9QZG0OUtBUH
EBBLI74O1QLHq9ohHolHRxc8k04wW2dJ3XaYT9vjC9z33515XxVcUN+vEw4u6y9q8FgiweLT5w44
Pk5aOuetooGEwg/4I1KdwJdjY+JokM7EcDXjDfDVjaDfvmhPWclEigZsBhAaFbHTnNiRN+5gmoSP
nVmvZm58P9dOiEQZRRCTkdYGnF8nqIH59/zoUZAw01L1+K0iMXt8vK7+sJd1Vtf/XmhGmrBJAH37
rSCrxFxtNT4QHEwHw1+kHHFnF/Yl3NlOQyGUk0hgwtJ0kRlnTIH1Dp5qTz6UsTjnBAK1jb3ITcXo
kcIogVrq2eyyiYdc46rwYA6sXJ9Kf44j4vN2SkPbn3+pwLrmjyYIh9Wu1HJBTkMJtRi1kJVNqwhD
sPXBw4AJcvNwCqJLRF+KQS6jcrRMvmiDtJJhJdCqAIBaOJwH4IKXsTEzmjp5mZEjcHMGRYW6TBYv
z27Dn2MVuC0V3klvMBEbGlPZbEjVS/XGRWCe+8ncbHpO2NKcurFXB7AVkP2sPvFd09vERNAwF7pL
i0cS2PFuaYh6ZfANndDd2p7mFpAi+/NS2oRItckF8q+94ITUjv6Ddi14FF111PIGNcURfcH45NQV
qmCtuACHuBscJTs02ZjkG/Ff4kOkBjJwHfN5pOuYnjUotxlkKjmC15m1kZUKi9EXK9cXh8E0L6zy
J5MKpaA71TZ+tJcJPcOd7+TM2S7Yi9lQXo2E6dAhsjp+U/dxd7wf5exfyLQcFaS+VDZCz1eQdc8q
S7OIzV1WmVUXiRID2Pefv03nIGqnLECyBLSYq0ns9YT3dG78apVJnDGAKSlD7U4Z7c4c40m+9Vtv
CeHM1YeVgAZCjSjrZexoN3CcvW+LSGkbS4STbLqGM1SfWef/rXNx7WWiSQthq10iVD2PwRTMyybc
8pjcxRsnyHpbnZtw/ZWEuzJR1kWZsOQHCdsdi5u1aA3py9IGHmlgFKzocAoxStoPUT4sbjn+nMUf
0jsLxAzI/MDzGqlzcd4j491CPDO+9056mPf34N8sO8qWkir62PnT2rzmn00PkkgRMB+pr7nlhPU3
9R+w9QlrqKwGv2cx7vCkAGB0h2gTHAT9E+MSh6d36oIQQfvzkllWKdk0bu4h5IAUjEClcvaaAy+h
ex5zFhO6a//zFZfivDwyzLX9gR4ANLdpC1o/y77nNmnlbpM9GtzpUxIo9SBh6IBUCk+k0H91+bu8
BXufipDYtRMg4ZDdwa61ubwnM0LaKfO9ercxW4AquCsc5yq07y9WAk1ovbg4Qvj16jStW52LKcps
sZgtA2h2qieIuNR76kLoUvEZqLHKsZfQqPwTyM775FcnQYYTHzHgFd5N9H9AZa7CF7aEdUdauawx
h3j2tJ1518kVYigjs/f9zphFwCK8iiu+oghP0JlMIlVmScZORWPtqeCCd7VcHqPl7dvkNTGYf1zv
71zRvXa60M0gYAeCOsGxqXq0wGjFPvPFTANwnAyqaD8MDkDtc95lLgapsFaiulSZupDS2ccDl7KZ
VreIg7V45K4AixUKfvMaPo2vQCqw9dfyVyk7XQOWBOXnSUV2uCTtwcU37c0BAjUQ9OuPHZiOpr+h
e6giUFRCyLzigIfayRWqBI6UQopx9+JYmpZ9j3hlrG6tK4ebD36z3aynj/bDemwn/QS/XW5Qnj7W
QA+oj/rJYDgHK6qNC2ZIFXbSnFgfCWhSP+jAlZrCjGXbOjrYBNBOvBNTC/kxI+s7mDIGR0tihP5h
BBreWLflGejPVt1a/MoPTuF2jByQsZKnVYrGUogfYnHXQIVtU2+IUc54zaFE4tZCecsbOEhdlb8E
xSdEEPIjk2oRB4NB13cKsweEOAtflQZdv8NMP8rMF4feHNYwmGmYimXDlPeXaTw4ioT13sFlD3/w
2MK9X+vWJe86SiYLS4EhW9x4/F7vVabCz4zSkv2yZ2jT777NCr4cCMyQSpY1v1aWXP9dYab8uRQX
rCjTQjxWNAc00UK9CmrFuml7/GYNJe1WCdoXqxVY2HXHWvyXY9KRZf6ocNsT3SEknU6i6g7QcrJR
22RHHBAGGlQa3FtLGywRjn2SvvOMdLoswh205nv6A60ho3O4sqgLdUohIFRCJdJv041dntYnRV3n
eSdyIXC5+9iJUQlGWQuXDE8/HMGBczaJyk5QsmAGtUOQwEpcw1lvIbyomh2jarNLZSIWqByqTzC4
AKhWZ0MEjtpJOlnJv2WqwgvMxxd5zh/PxOiwS/EjLrdjcP2NFsiZA08g655QaiU+fvvqhnqcDFwJ
qf15PGVHtwEjvK0c4eNgbT9KhOJ5p/AbRUZXL3EcSG9gd56SlscHNhuF68VsGloRrDHMDfZqu7NR
MOv3scPlkXXo1xENS5h6mUA1nHN1RNmFADNzQumbW0GVJ3locezHAfP9ZoiAKm/3Ms5+NwWzJTo7
tflj7Om7j2TbMOWtaE6Dl5CwCJWkDL4+/q0gqkmQ1BpMDfsv+OYyQPG3J6PPa0mFX6Gc3A5Sas9c
KATPscPCLz74OFnTc/T5TkTC2T45pPRgjRqAZthy/MSRGxzY/mWmz40BvomkIPA9eNzsZWxOfHc/
Um7evgbLO9tsvziWmo2Y4U8BvRfhvDh+cUFsbMB4ikoMtv48AjJQBrTm0FaxpEKhz644Es/x+zZ8
VxuTpIBvZ/IjTxlDfznu1edAP7egyDjBrrPsFmdIRby753d2T2pKEj1l+3wNPa/N42/ZO9FedBKz
ft3R01XAYnjiBwFQRNL+Fm7o2Ojyw7QVmXEWWKMDKb4n8rYjG4aR29D02Rb6XjwQxI2iIhsbPTMI
4e6JMqo8gs+GUBmhln96tmSeaYaCYgwvHWJYDHFNul/t0tj4hn3/wOMftUHjuaekLyyofeKQPcVv
XReow1IsPB/x/9d2qtPwpn6tfev2cs9LM5IKpK3Q5YpC57qD0YC483cqRtiaWXKb9WjpGq4QOzqO
DT/NWhTaYwXzhUgDbg1rSNcUfaZj0mUKqYd98PUCh9qe4gZdmqpLW3VyDT+Ez4SZd18ufxb1TWQL
5SQwA86IFrXxBPMbfK9TB7wqS8L9COVMhJUjlvJvNCWkG69SEUwcmFf1gflCpJ+F+v48GglfHXLR
BcHPMivwbFW5OwAs2i91Sfff/RdUIZm7v3ANyojpBQ06YFQCuzwqf52U743EONIwfRL68F4/2uVg
zgXGqg4Xae1EWjHic7MeWlIWakpxL9Lzrwex+AmyuRw3w7d6y68qgDQ5tA43M73dGvZIeexub0C9
I69PKbI60w4K8Ih1BnxIP5KMqh7q4QDJRIpzNJGowD8912BvQ+HrAa4CM2cNkw4btMQExMlgEbqt
calG7YWKebwM8UY3n8W28I0XZGIuZuOLf3/dokfTp/z6c0ZPl7XgBKh1Ieeuu/nE2EFxKhnzR0je
ejHl8PVEMQ6OBAJioQhJueThOWkfPaqHevQG4Oa230G4KNRRhNss/Av7D5UxmltPqiGcdNVNDodb
Ztd11GPCp8jqEXe+Uj2h/fkkzRUE0GlGgrfBMDbe6L0sVy0jw7E17bKEDlvbgJr5sd8nkDpKMGEK
J0k0aU6vdjLjDeDhMlD5E2A+jvEee5HTn1CpS/gI4KuSdUblAH2xFmx2fdK6U/rzeWUoQR0R/Ra6
4vXLmFhKgPsZ4jYptY15dzqhVl7idsxNT+9G19W41EN9EZwlsxpfJxhXRx+M1cSj1HDNjgE+gJ5a
lDHyW7IKgn0sNlG8581W1+96LrNkNkWDIiotI+uGmKQz9rrOt0JPn+hz9M4w2kQaPVh8n5S4gnZk
MB1I8J42ifbHiBG6f/e/jIOyr5VsQB4hA3Rr6o1911zdVorXGj8OBRLXAUjL5YRwpsSruoRUnqdg
naKBEmEfgTSWweDFWiK8SBIZLiUNOIiFJbnr3xOszuHYZibX005sxD8hPlOGk9dGkKYbK1S2fjEL
+4tbLjTEx6wHXyOVlIPSvey8vx3DvMKWlYElOcGAP0xJI7naMgcUGztVH+hBT5YSJGGFzntFK1kf
GppuCMe2EykktyquSxe/kQuYoftf0w24ev7a2WadA3jLfskfHtXd8X6RxFDhRL6VKRi34FVMIP+n
vyvMXDjGmhuNR1GjmMEFF8yHl7vo+u2wfdcNhnt8NUrlXLHZ0kawnOPNm7hM+5la6SmRBsOCObfQ
SUL44iKRBfhAF+GMXc/H7fHvNSybAbBRxr6el4zr28Kebiz0oqXpv4SrRQJ50rpfbZeRKhu53XKc
x3pJNyP9rOknGeE//teCatfQPViYAhZMDZgT39H+u2TJi2xF2+zhLVgenOy3fjdzesFD0CgOEICb
ys+JrlqbTvt7r2TX6ChTfWFKLBHuUiBHuvIaodFqFmZbFv1cQz9oKeO5duJpTkxCt7VZsYkXt03f
SQxluqVyuZzqB+ksX4zID9Ylhn9m3hVnY+NexlzyClJXkt0OGfO40Pit5SO5MApEypcbuIqmP6f/
gaYjmQbWEfrhvqR1/y1lPniRyR5V2fdHmhGdf2DU96ZmFVV46yzqanSFMgXMHRSsIFSD8BOhf7Qy
dQg6M7yB8nLglqM7VwsPjYJum+Lob9mTZE3VNbhN7UH+7mNaSbrPnWPiXDydxNlpPf7HZOraI/z5
qdi2O6yj09XXqrBN83lpn8q1bPntUWiFYPRO6e9NomfaXxsacN5lAJn2toH0oIT+z8DzQcs0Mld2
xQg8jbzmVnr+IsajE81Z5Ejz4yw0l6T/R6xJLadzUc3WL2TQXs3Ur+nH2+MpJ8B0zRzrlVhC+ozM
Ll4vNXj3HHeG0ko/SkPwJkMX2anlunBi3e+9dvRQIS5el0FJk1+UbWqhbaH2MnygORF304caAxdS
RBkaFtY61ka86YeZYzJpbt54shyAHgX6xgQ988z0VvMrThzBGkzmuZ3pb8+4yLny0kPWyLyUWPgw
UzrF4gKqaP2GrvI8fLnu+uG3ZcHGDjSo/KpDT0V9RFqqwNUZ+lJn/uaYAfy6zBuKGKpISHfBh8KX
/bEDaNrQ2S9Q6OK4wJc+L60+kvjDqZVWLOn/+lxgPFuuYuu0oyie1Z8S292lO50GjBUDAV1An/z0
vbkPiNR/W7Rmu7wBmwV+8pkdmNEpxw3WYNfYimp/oj6wssPNU1JjFMFgYAXnbWrgKqTmr/ni6ppY
r+tPBAYHWG/nPODJYDXcNjJjMV/aKDeF7soAc8CwkLSbT/wtuKD9I1KDp2iynhGpzEtUse5QLalI
QTO8pticjJwVosPVvijKy4kBBvzbvHXQxMlDq6EV1ly/IAxu5NWSHxUO6ykQyISb42WNj435fjVr
NAc/5Cb9X0usWsK9QJZhg1pQk0VVk5yFDjowXU9HmaqtKsKUvBTDLbrHx42RvxLO6BGNsnT4hGQI
1ookB3L5vPDew0APCZ8FOhDd7MJDyTfEn2YAL3mUbAEdsolIuHZ5GFnhN+xvkbzXqcla6BqGVerO
IPO8gHFBu0dsaWH4h03ofA20D1XDk/2h/CSdvltUvrRrxb1iwxuN3qZlQjtxs5Rk1qSfId+0aNTq
ncUO0gMlfPai0S9diGK4MWZeFUvYC/SCjHpPa9h8zmhsyNohGfUN3LM29JLL9fN5s+plxMFvOlo3
HAln7HO9H8Yf7sB5sqVZ/KjbzxiCJ+QitHiyARK8SH+xnWMDg70se718KgoJ2dQ9dRmaz5Mu7AJh
AcqVJwno3FmPFlwEeRB6EqiLoSur3+g3fw/vTYrb7g280OQnRE6PgOYsBd8Au4EYdp399ajjxRtX
q+oL5S39Ewxh5bOjNGlx55up1E7vIDqfIptT1naheDnaUpUejahKsU49LXvm+KrnCJ94AVjmJTN6
bqQuu3oaBRl2edwZbyhlo93oaU4CFDfHOT1E/9oGNZlAPqSfPCKPxpvct32iuUPZw+QgvaDfEvTz
FXckwhuL1YdV9ny2yTnE/dtzu1sZin3PQ6C8FbPIbUFRqv/3vsWkUuMQBMF/6XyBmCkXQoCOTB1/
AQA35+W9JI8jbbRETf7///yAGS6CEZSdv+BfXn2eZq0xJxc8TkT+/9vVeBqB1wWyXMyeqA3zcCad
PPxDPv5hNA+Q2+23JWMPFC5EUwjjgLzpJ2aZrHHYjINS17cGVyN2KqYQRkhYYgrPzVo0FTE34ox2
7XDojRInj4eDP8ZaT3LeyK8NIsn54nwXzAnfTA+32i/dtT7EVjEcvJjXg5AHsRufhlQUrea7xBPN
Psp3zgs0kDFt+DQG3scBufPSCm5MB3EVU+rGiUNk0wIBP56UAQ2Nyp6qHFY5cB6asiba4TVAe+HN
4KkcO7VbauEny/9t6gQVwFjNdyOSwPhN38dIBvbS7HDkCR3n12EH7emuXeZbP5764HiUzIXaJ81U
SQnaTQJjBW0dl9YpiLviymAtN1x6Iv9RgBEbWVFj0vefrfbvEX3W/ab5DFdn63OJzgpbqcx0VKmq
ZCN4V1i3+wTFf/JKLIajn1sDNVq7Px/veW/MmVA7Sq+OYk+LNGHjO4qqzq7T53xU4z8hAjHzzqHM
eoBgEXv9pFZANKtXIsOt77ddlZXNkAQ7hK/enGPfyVDfOrbuJiRtE5pky+glmWLN9Jdjb03GbD0J
3i0ZArzbumxbrWmRcx9QT1eOcmn6uP9R49T7aADIHl3w+t+uhhDrfYszfR3toL3615KVz9vDYbVM
ksPHUjiLih8Kl5r3rKnDiOWAiM89OfHUBJc0VeYDVcy8QS7d8zmJzR6v/ehW9nTQMwupMiXHi3W4
Xun04qDp/ntRIpKM3YUXZk0k4kQ9pj4erw+/9YoNxBYbfKnWsZ95rqNonOWuEwFfhW1reSPaHH4l
Ea3b4A4xaEISkjfE+dNaTbqbUkvKLeQj7j+6HF68SElukCWjGSqMleG/TJ7lRYti3kAAvJbJtuos
OwR7Xc8EFIn0Py717xiQfxsG4OQMy13BEO+h7D5IlMeW8+vUqnrmY98rjs6tVeoaeqsku9fEbu1u
BRot1qGw9DLYO5/jUAoBCCWPEBOtn8BOAVhtgjOlX9jEdVlu3raL+RVPKctGXMvC49OYIftCEIE+
38lUUqqAlwZcLPpebL19+dOfBco91r/VsH60ms+tPuSCleTlgqUzpBc2T7YBKJMkdgyKRjIs3Vbi
onCK2DeuceDk+/hdvKPLbDW7BPhbxWz9dUVyQbsK/QTlxAhaBYJvIsMOdCmUd+IFH5RZesaIv6Dq
yESqiayWegifRQl+byeUWEUzPXBoXQgzGHBDK/53JFB0Cex5sfYGoJYdf8SgXmpSGWGom1i9rGwS
CS5ntA/AP1OU/xn/NdVBQ2tmYgI6fJ5nmZrNPWYIQLoi07C+JKIfWjbblyvs46ESQtjZAbfvTILr
J4T8Gu1M7o0HE5DExTj9t2BPhNtfxZuztPoaRu1F+t9zcodSYDEKhy7h6b2eEi56541IFGYox8Nq
rN/dZU//JLuge8vbAUVxZ4eXb+382yseXDDnH4k6nHiIDC+p86jOtsXyD9Lp7KDku8Chr3PgpAqY
s7Qs9Xf4eKdSVUlTkWfNRLf5lpk3YjFfnVJ/JMLKSn98p+czWNLOO3JN1fbOk06CSg+obQ1Qf5VR
5dJTiLYuj1+Jfo1m5uQBPEnP0xSiWVJPhkMK/eUeBnhiGtvsGH0EssVYEPm81Sv8Lou4xIynT38E
UBkwd4KxGecNROfWPDoIC3hGLWZs1ZGnwPWu+hkxLFJav7wFAZW+qSRTCKbL7FSg0LhEQiMWlZYG
D8mX3CUk7Wpduohof7fV5WtBZomeiN/XbmF8Uz0kXOCwsfrG4zBrHvNpdam93O6uwcK6MlfCBykn
qvkdvxzR2WPHnNYtPx7scoOpV70vagxHJyg1kFDQObFBqABG8cksTtR+fiSvqS6j2AErB1JA2QqB
Hsglmr/T04sRlcWD7ki9T29g6Kn4EAFNRl2qYiyplY+WIAI/AQp1tGjwdjOxdRxEl1rVkLfuWb7Z
vRICJfPrQRl1JAmoBcuhKNKfEKagpLvsPSWigLJI6V1sMIbdXXZBAqJcIxVZkWMXpZAu+U0V2Yqe
HSv3IYIuSbJ+4RNJCd8IE/mjzGELGtRDeUkeBdgkMroK3mJr8Vv1GA7DVLMHLk/YpyR5XFPWjLn8
U9erXy0EbeU+zZlYua3jVFMUM3JQk3n4Ovq6wCrOVLMI+EINiml1rC2zKlZwacASH+W2fD1F3Jei
naQDsJZ3bsoQBQIPqih6q0+yKH94v2t0tPkaUl8tO34BjTzXRrVAXeHaLUzNFQZVaKM8f/UjLchA
9U0z23qbY9k/C/XxUv8pdj7m973m/bzoAN6he0qb00KOTopT+zR/8qY6UcXQN00KGXEO45H8KCzH
gC3HjQdUu0j6fLcLOpR66IFFfgSgTf6FY68yWs2n3+NzTEEE4TE22N3rmq/wWFeRRFoTfFxlGBK3
cdAnDESYnWLyGTVy08uTxg6d6Mr3f16N7rrVv2rZtP5OEuznpZbdpZ9vANH1fFtdv5tibbwhN2ro
SQAMNKP1pUrUqIVZMoo+YpVXbja0hoYa8GwwmpsHz+snFUgteXE+AZ0XE3QR9IHNcgMnuAZ3eP5o
Rqu0+ylqZe3TWaOyDlAmhKHW9iblWTUgKHdw8bgtPgLP2Y8NeuDukItNBw4D/s3mrZY5xzgCzcJ/
FI/5JxxXZoLy/jnoLdmZHZasrbMRKGNZVdSutHjViOd2GVCf6TtsQ16UenfhIDGpxlnMemhF0OLO
gsk0Rhl0690YHIaLluJoWnH8uEl4F68O09R8y5FP6kjY5OpzmxGK7ERW8n4yJ1zxiUxx4o2/tWtU
aipfkgtcu9A9k8D3bPDDRLmuc1m1pMz8D1xhmUn3QdXD8FaDjVsHVr6oz+9t9kJ279plr17kBTdI
bf79/ymjY+24PM/VzkmDMoEH+Sx7SqhaHBHOmi6s0oK+gcJAEKD88iy2ks9vlpX6e/9bRupSB1B4
K3x//+yWhMg2A/DCD/HkA24QPlx6JWuOvxoLFT72LFdVpFWWUas4FszQH6pjXSybNsBn/OtUdrV6
1mmAaUEnWSpfU/0v/mXcMGrQZbxHENNeY6uQiYG+zVEtuWvY3VdaoqMv2JOLSlEY/YJCQG3w1VqW
ra5eoXznrycBCDxZ/wUeCmtf5ESqFpp6xSLqVLn8b3Zgsc1h2DTF+20RG/d7OUz1ifrWTsj2T3iy
rJOraKPkSW5+gBNulCZOSnYdFcPe8EIn6RMkDeWzle0fNK9oqiBaCTSKpuFlyIfkUHUuhN1ru9m3
Ds0aDeUpCu2yfgwwq80P9U+pYzdue3md+PgFTGfSijfHoNSJ6WfpoBL/T3MIJT5l8s0bnGW7FEAT
Fa264dL5bpcK7z38tcPzbvC9y+R+P1rsIlRSxASUiP7+iRQmcIL9e09vhAajuU/ezPvoD/lzo8x6
bdJdyM9R9MT1F6scvJc3kZ5kueyFdDyNoTdIsrTpkTvX7KmRW626piseX/Cv5PxzHO4Khi2lWeaS
3Licvh/cI6o1OKBbZb8QqUV6Qy9ZdEh2H1uQClUsMk480QqaOG7t+cilUClSjN/mZ65UiqSk3y02
I3M5Ol0SToFEsoTDZjllb8gQ8RwIds7kIr3Af2etSdhDqcDB0YiwlbMz+gAA2gAiDo9BtaI99Qd1
iq/4D7VrIk1wb/RAh/1mmqZ6menL8UsqS+IHXovw+RlaOVN6ZK3D/He4VgdJC0b61BQU+jeueYyp
KInSzMiO5wUoIecov6ZfCbjqTlGlZtzjOYd6E2WD8H0+PFrJooMyJsA9et9SkhnzA9J1pRute3Ol
7pEmO0SL1H31/aoPiHSkAc31qxKjOBBxYiaQHAA6jj8jv7VcFFR2QBKNI0IS/adXf7BPVVJ7kA6m
KyOzi7kZcSNXwyatQuxGF6TJpzC+tlEtnecWUtDONvz/eZrg6PCT0/dOiBgGnOkaui/K+DN0CD1F
Sw+StAMfUnYC0PbthRQEUEYDLNft7XnJ7obASuczygjZPQ78ZvIXDyEfZW6TqvWp+dbWk4pw0kII
FWNhhRgBnRmeTm0ZgixLrGmYtNkfIoHY47FwnXxkPfoF2J95kH4GTLoUi9g1hOijMftk4ZqV35YG
bvHWoGQkubjVW3d+QfJ9UKg9klKVJ4cLqYF9sFfVkl1FjiSejFGvNC5wNyA7H77Z6Vz1d0+oPhmg
7R7bSHWIwZxiQaELj3tY8m1DPhxOXTKKKitCascbf5wdX6DN6yVXqWzXYKWt8k/vtm/VVxu9AH2U
42ozby+3R4FJ+gT1kGQgWA7TGYIsCKoicklkZmHN/KcBWRKfLdmkPMQJ3EdppIN1+isqjmpAwBt9
wV1t7Lw/Vbyr1lZcoUSVYN0lt4ZJ9wGu51Dz1NZ6KgcCoE+7KB487XbjkOzk0nWq+DSZgA4CuSMa
B1MiEuqiO9r/tHl3m8uYEBKArMw7m3N/rbUNdoO4bYyIdOcPQm9ECphVSQQGrMi/PWHwt0KuiGDu
4aMZAqvRIqjYgJSSfmjZEbyOy1T6rRs1G57YK4bZeb4lkjJcF1kbDYx5pBn0D6tmG4XV5JCe7BqP
0+MwxuCFUdyklXafzMVYHWKrCkvSNwRHBjeyXXgF7QajsVdjkCJ+5njnGI4YIseUx7NHua4vqce+
QDij9kkh1tLisacXM1t8YXYu3YnCOU8h21q1KgIPF1OwtQowMZjNOkpckSZmxzxglNdfMxY2Whc5
a5vqbqgpJMhFnzwlFyIdQoWo7dD2zhx87lEPXHn+is9RIhcz4Uj6w1Qul2uHhbWLyS2Kgh/CxfKr
5kE/q49aR++9w3aY2E0qG7waZ0PntDfMk3FYJlq3MwZFtNTLxCIIMC9g/7Zc1fke5ST6i6U6kB4T
YkJEq7cwcX0BvrcirtlYcLFV1i6mVBFj85403XHodsCta+jIIAi4jStQSqd5lL/qMnfRLEmr0ENd
elv4Zrw/VAl5ZXAN69XwSbKMw6FkJILImMFXO8XQLtQTwpWhh6DUMXxGd/wM1MtcyuJ0/J36+ov/
Rf991tXddu7PcTYhlAalsZwSGgvU0PUA2ozmZjIuQ+gjVfQKT5KOy7cOVAHiODt6d1uyy/cyewKL
0Nb8/v+BkNE4hnkRGUV13BHbAlvA4/BCpiLSaO4FJh9TOTZn31GNMQ6HxGNSo2lZrcGHBIz5VvDj
KYGnsQayp/niEwE9xGgHoMxKHsuE8GD5gwaEFQr7BAs8yMOw8MMSpo/7zYSra1V6KDW0mHNvv0zC
2/+4SFtjQw7zolO14CoJ7IwBYN/GGzTUgGm4/5ng5cXZk2vcSKftt8cLMPzr09jdmkpq4TvUIvWp
svn0uKThtiPeZynRm7LOdMKMAl9T5XPHIy1g1QMq+0j0Weqmdm43Z2hHYea4KJIHCHMQP2oGFRpZ
WbUYGJAWCOHt/ytcRd2MK+XBfv0Eqc/Om/293O6uHu4XpcMy2TdZiMy2+/KoTr0eZrXDDtBfl5t1
KvZtkO0FsY4ld/ltFySmQwvPhCm9CjXcFH+0l8Q/fVRjvtWNxNCuunTw6qu/z6PkKQNZGdRD5P0w
ZBovv3XFaGmAuJmG1pF3KETgdw5uIeAKBkoje85Kr1baYviKrt1z1kRu//QqTSaQuzeUzqSCW26k
gZbOma8Dd1k6rgpVIILFBZAbL0rQBdIFF/yuVujSbMiD2wrDhbPIe2YKVUxS74nxi+gmadOPFpcA
Faa6sZEyYl9HDo+mTdnQ9hKTnG8JOXB7XjHlD/6OcYLamPQdACdK2RJNpx/HJtne6CcGnlLgLW0S
RYhW3ClBXBlDms3psxeJ8lce2sSGXT0R3EbNklzSLkn5mDpHwzL50S70DQ48cwsRaF7KJXCOK83K
nvoP65cNOlgY/twtw2DpKACu+a1w7GC1nOrgfPBMkSvymJCRunXebGBh+CJ9ExRyMnYv8nOzAMiW
3zT/YUmPP81ChnR6PnDT9uF5SPXPsuWhL/hiORWzD+razUAf6vMlYp1LnIewV8zTCJ8UpigLHsAE
xfnjL7DN5ctQlpVUTbYgTcLG0bu9Nb6vEFN3ELAcYOLNZKaNVVqDWcdnSQzoi92XVBL7x1WP/TQJ
Viq8J1Ckgpkeclz9JAWmHj0/m16pe3n7oHPmrNK700Alk7CjtJpPR2USCB0aItv3dpRhzR153y1X
J36BgKGvKuhsBYKhC7UUmGvAlyn6i1yz2RMCpUovlKrDigz/fACT7frkwM/QWFY28tryC1DHcQwl
37m6HdhQ6Jka7kI8BJtivZvjoYT+ASRX8LRKfKFvlLgKcd5p0BiN3vdpWlfeIe/xQy96QUfGfksR
M6vW6qOBPzUokrNxX7z3dUK7Pbw9fYyilbZYA1UlOYychqhnFaBpv/WrZaH/SEKBOxzUKHxDXalo
CBzdCpyPuHNHRZSmKFC5yaBGOYt77Jzoz29jkJoJkR5S6VzHvrHvogF7lE9vOsf+BfCTD6QrpYrV
F4K+VkuPvQMV5eyC8VWcoalZHWVnN37AZ9CGSW710XSM4Yl1uL28qNorwMoIaOeSl96QsOZ+Iq8V
SgXtUfAQTcqvmgchkcHKZADEmcQwUApD2YHEnhzajtA3vo4qX6EW68MI5VscEnUYEUM5BEK+hvqa
cNzJyqVloPeiO0VIdnmBZUTMiWWpWfg3IgefRhVNlejKlV/ZU+gVjHNuVXNG4RgFYB3aOpsHJWTN
NpvcNbl0Uncko6Y56wFyY2Xp4oqsk+jSDE9mDNw4NVrcTGCAwm/C9fpAr3KluADcERjqYcTgoWf8
EmY8K8ZcDSJiqaxIXTjp4EbhemIwLA/9sJgObqTbSCKqZDz2GmxGNPI1e60bsFiXKQ+Ubt34omuk
79gOBBUR8NvIdnN1FPYv865ZGrfZ23q33V14mQz/BksdhLutMXveWPYrB8YqJAtZ0l00XTUB3+Q0
g7V9R4M28ka7Br4Eckh9jGIX0zs1k6X/Q0S2ChWuqC5Z11er0owsJPKBOPv97mqELBXKnysojliE
vYi5W/0BJq99uqKwRhI5pzyOq5kKLoDRzst0jY0uj79y6ZKOuFqs3DLFwJ/5/vpYBoRzm6I2q/lZ
MbPlawOK65TZKxsA/JdzrVEIR1uqGQ5u4LXo3W+QAEZC+kVsyDmRsAm+COK6krsG/rnBjx25BuUT
mQO202JE8MIY1UlIQzUU8AIZoqPe0xOm+yH6ngXwv2W4SJFcwqqYBpqdqEATUVrBXClJ6uKW60CO
9kG/Iiv2xOXTXxv+3AR8Yh6n/w6ChQD9jlthQtrq5G8w/qA448QnAnmNfZF7xkrZE3FQwvUOkahf
Kdb0UZG7YckrcgQwr79le1fA5q+OmGvVcFk2m0fgbbZDz+B2ei8PGVEwcYTBgBs6HGYhWhJSa0Vv
6rB+Ra2bkiCsJWgJnjPLkSr8vqrny+cwBOeKnaV58U1ESF2Jntm98w4aOD4LVzzLAUpE3KQ2kfyA
GduKK4TvQRprQH7YlAtvcD3mRp6INZbaOA0xXtWfHS2ModVmpPXSSs+SZVQlI5LDgzQ1ORDoJvm8
8pxCGuF3PMzvhRNHGo+tKjc+E2l7dG3owGAUYVlUuwyG0S+dBrtvH4KbguydV0XnAVhlVHeMlfUK
WzwCu4tVTGX3Ok3mCIESNP4Yt5RrV8tsI8//Qt87DFcgrIGOPoAs4smMCEQ6xGRCzzUyMS9iRBnb
TECJJ66xdyo5QUtKd7ZUSzhQLCQAtqF+p5HsxBo9sd0QYJElV3+Qa3rRkvndMePptLTFm9q1cU7J
lNrq8x6d15mnpb3gzcHCSCAiI2fk4cJcreqGDrwTMIAoaUjzyWoGN2dJyelXk722gI/5y8sWfcsl
bGYBhZVfFSz+GXZMthzk2FtpxteBsxJnTpT+IPPZexLmglWdgoY3ASgi6FWuUICnzs0DgUGnI/XJ
MUGT9dQtL15ZpmxL58M7vaUIIH4Kao7nLZKeSoIgrn7BKs0y/0uW2uvWgMWPoqeaCPl6UMT15CZr
F2VmrdMaCklnfSbputERvGM0cQxceMJ6JuxBgzKZE9Z5i2qMivmPKyGE5nt2CnocqfEO2/gQB6pC
JVvOuI5AsOzeJkAA1ZFMvHwkbEGMPbNGuBWBmYYKT+tiT/Kyry2Pi1ZuPJ1OwBqwBvPDeHnH38+l
AGL3wAGp8x7xL37BI69zA155XWF4ni71lnoRpyFy8hoeRJYzw2ohrvlAZOM01FteYpAJr5VGlUQ3
B6tTMJtcZx1GCu6A7jXaCc4RT2P9+hUn2x8ogcE6lZKJgTkJBBV2FjJahn/pnYlUJjv7PT3tKG8y
+utHLavS9BARnCxQLqCAKlm7yBGc2iHUcZYcvtUkF3YNxuVIIi3YXiygHmZKWJoh1YGW7Mc3hBMn
2educu1G+AFAUhvOTTew1x8PxiR1LqlrjoyFx2LiSuhhlEU5QMhj82NWV26ra4KTsIUlbBOaQv9u
VsIfCFcsccymA2Kiq+SepVRqyVPeAmOA1fTTKP0iN6sHoQXVKtNIdoLK+sTFnezOEcILSC732+0M
TMnun1n+q6K0tPsvgFFZy1ym8atd0+iAbGteykVOlTJkIzl/wg7bx/rAHBagpN5Z5ZRhKAI5bN2s
FHvmPtbc1v2I4y410SLljaYS/5xjLI9SG8Yx2LqqZBsDabO0oKkKuA6fBK6jQ7ZD0g5PTFmmrc7V
YcT6bqGuOe+b5oeWcIa40YLLlBp3tzmHcTIKBL152lBG9WAR1yeJV7BQWYSg4Qdk+sWgChGg91Ca
wdg/7AF1Uom+E+U08fJgfxgmVWptgDikq/6vTGnCLsRdTvViuG72/wDWIf7XIj5//usqothRdu1l
eBtF41q2EAsUgBVQDUjUL9qjK1y7mRJ8k0rczYJ6qwSzUXdd1W+Zu94z1DRQwNjDocZtAEQmSnoQ
6iewoiABpRGIFTlXtoOaUmMnpBSIdMxIEqOl7DFRmPAASpLHUMaAQ3HzBZ6g6lJLBNtyh5XuRsMu
2IpVYkcGewI/SJQf01FrcqAfnKCzN7grF2wEBrEZKZ8ihhn06c2qk41PBOhPKonK+weDv6bt77IE
0XcLVySD8Ar4BuskAlZliJDeoaWdfj7vnImOMi6AEJ2OpOCy85fCAxfnvmweIYOah/jNF/ThFY25
L1jAUlFXekPCNVVZMP32iFlhssWzXz4N8AwgdyDSElhcnfn1jqX8hvp9zt2MKJ/ExCI6iR6oGiOX
gpFqdjqUKU+3CsmtHTmj1bnUBImQSv1G8TdItpKVixhJZ2lDk0FP4+cB59Z5a6e5Wjg92q4cd+kL
Zx53rEh46ctArGnxF2g2SuzGGY9fg8Ev5+lhiGxaSYV7pqIOgomi17TyynsfnrzzAWcB3JbFnDVA
9H8V2qBR1SEpVEja504EP9bsjIyJQII6zCuZPg2dcVLiF7Rf+T2Nay+6+7MAVenYNPg3dpO/EkbY
RRdzabDsrON73tRdDHlivCvQEDwS7uD85YBcfvCPo2sNYWTcaB9paqHGCsJNyma1y60qwHyjclcA
RqjjTPYhkk1/2na35VmcMVxSElaW1tipLbQiiOyIFWH2F9LrPvWq28FYlPMOVe66aN+6Gi5s+coc
Tq3RwVYK0YOMq2Jm6sb8P1mH0xnUPt/g/ZITmxDAL2OK5lmGq8N/qa73yO2540+nPe+wSBxB3his
27I8sD+ygHxr6o9cnq+2/SKlOjuwZLZbEqP+qrWw9vk8LrDPLrFOLViPj69TcLFGcLSi7m/4VllF
P4MMb+0qMQHOPUOK6/Bsr3fIoc/7q/Dn5tjzVoXqpsbXcxKgQ9p+PkuPUpnZaxKuDigtG+VsfYDk
WjAtpMuFH6zBpVYbeyDv1/nAjFKh1k/7PJVIW1RjyLcnvfIkAgOxrUOaI+3DLDvWIP3hM9VEydXH
nLI6DlcYYuWc7K5lvMzK8pdWtS7WYdhgZkhc5nVfiKAcLBotwfQXWIstRpnWtrCCt0L1rMOOYD/8
X5d0TrVwvkRzGeoKCVxGzSNmqUfr6ErR1JESjYPcnkLLKQM5ZYgNYvYkDwKG3bSHsVooGSsWTSLu
wzaAN4nXiPwFkupUS6ukjXApbtP0HinvasruAq95y1fmq9vY+/qpEm/1WV0nXbJtrrWP2CMKNyYO
k7ILdoKHkj4zEbVtK829UjBBgi7Nbgq5DQ1IRrFTFAgk9+7kkeLTRmrG5+gemUlltsJK8NbXTEIG
oLc6fz+eQgnz4Bzqn0D5QoUIUBvxw2vYwEI7Cmc4OF2/iOOhkBr2nc3zAbFgYf78NiRaJcjR2QfS
zjA8XcioyzOzlBOFaHtqw8k/kYgZ9fGQi+pzuoOZTOd7oU+TIm2FEVpvk5fKCkBLcX+hUV7htteE
hfhsfru2hsuwqH5NsOOoK4Ex+FSXP7xIfuLMnFNGDflLMM073X9hIwmqyxwuItwWc3m79V7Z8aWT
288FiqePuBZrFNpRfNEyrBK91SbUTfPXDSUeSr4cEi5WRtjsNU3K95p6oIMCwv8TCqK8vPiAGEcT
C/xhdAY8wE4HU4GArfFBMf/Oz7bpk2qlOOkJP3a3Of51iPGZF0nSoV9yErFpDL8uzhJ4tYcwyl/y
TAEAsSnW2z7v9s/P7tpl0dqB2LVG/3z8Cnww6LQUaPWtzDsD/I5uqoADsdPGG9fwx4P23EVpVzDF
DNt0tHomjo5JgEBISdGYPktqtG/dp0Js1kPyeKdUUnii+PuqE+PBGp8rqu5W9cGhJMchpMzewhoO
mYYqtOLQbGaOicCmSFxVgSga1uRcs0eTt8K5k3Wk4XvHjQWSSrSMeLGAZekqfDEp17S0OYwamEIo
UItl+Q2nncxRHq6ONbdmLgJdmIE6h8tV2m2clsbqep4XS7YWpuqxnRjL95VUAQJs/ElZ2lHYRq4u
fzqcxaBTary++VWqalefF4XLj3z7ce25gRKFusmaYIp7m8/5DbAxu70Z/6qLEk4Kls/MLEZFASOi
0vWoDU1tP5pC4hGiPrAoMopfoUrDinw1lGbhrQDFi6E8gn53WpM29o6U6m4F3xqz+B3K3jAzgYgt
Da9sD99HfxXQfOPAaKGCVt+N3crLPVNFcyWHp8Dn3GvlikhwB7ygVYd/zB5QLMkoWiQxh6DGgLvw
5cASBfL83/HYZ2tRPrdnsHc2zop8QTHP7rZKbDhBBYAygCDBTVque3n9WUqLEtZPnTbU7FlUGtDJ
ucelqrRN0mxTlMocZsPFamHKxFYwd2CPT2RO06+jdahEi9wAVPUpPs+86pgwJUZIIH6NMKBlgBTS
7X353pE1Ci7lX9j3ZUbZ/mHUtB+cDrgYHv+2ieem9TtZJfgDGixASvuhQfcW6hyIWkNl0ilo1gNH
58+lg2WQEI4/u9HwwfGbfdM+mFnVyQcc7YkaqKwigwHPMvDgWKlEP4Mdlox3hNS23BMVDAdb4MtL
ZYV5kLILld869PS0ukoMb9S4FJfYXMh74M1JHpLsHDdzIRfMvIzGkENFQRR2ZYVe+5jw33tlifyQ
NByDhPO2jQoxjisb7LjpBwyj6uznOkocq8lMLA8sNL1/nn7Mvb5DilSaMvmgycoEVIT47RMN861D
gSeuKDsnyIuBFK1G5IZt5wz6DuVMp7Ef1E20CD2rRmtPZTcMOUSAmtgMBqACCftgrqCwJko5xFlr
PpUvvDWfB7nH1ULD0t77u+cAZbUYOwgaonyV6fnmha1ebWPcuAUwZFVE0HayXW9+Qspv3sdosITm
vK/WlSfEm6+odMbl2v5wPM28Rk33DI9bW8XzvqIrtW53XJNZsWg7nHmQmjHNAvMh+Duog98moDX/
RBnqY5ceRLoM9Vv6kA09wgXBNaro+Dir0ZTLZblBcaySFoXIIRUAroLEl0WOPDglNyr/Fc5j/aGA
A8YsRTzeaDlAuCj/4sZiOAaXT/Zvc2wjrv5nOVBXBtSAbl73IJr8GhKT8Khp+YYjZ4JreN2+9B2f
CpeGYLjGbAowJMKyyIH8UdRq4sLV6PL9Ed+ugqevLki46v0XQDkInt/1gUfhMuQfcs3CmakXNcS8
kxxQ0nOWKBxpZeL6UGsbn4CR5mNbUkwPaYa/NuuMfLbTgmnwl+dj6DieHu9Qpx1eKM/aI9MMzUMm
ZN145Ct4b1ad2ngSpkXJtgljZH1yNST/jMFIiAqpLeeF15sOX6fbTE8dA6KSQN7OLSxRIdrdcEYm
6EMBTnTmgQqA3Ee2bC4XeNkrKGjcgmCtTwUEoPEcbvD0IcHQE2MuS9fjldDAIH5HNEc+vYGYauHE
Tcoa8wz8jLd0sGPR0snS+fMVq+cpAeXJD290s5lc7jfOae2E80P9TU2gnf4h17WB5Zz5J/V0X8hV
Ku7Thgu6os+nDnLmYa+rhhHTKvQN6BCoSRN0iAj0OWGo0MBWrK1kZ4thkkqZslE/rJe/ZEmU420V
BVGaEPvUL1LLMpxIS9KsGFWrkdHVr7ymzMRREbeawAz3k9Zu/Dq7+l/P+H4wV6KKGos/tRFfeZ18
Mwst1KJiLCtsFOxCAcOnegM+My2aBQrpBjWer8OPhMU9Qj33IqtvfiQZNr2U8cZTRh1mtMn3XvNj
0pvs5unU+EgMb+ksZP4nnkvECiQ0G7U7HvigHMKy8rGXW53NFRGt8MxqRsJRmMmN3x7svJI7yD8O
tfP3zLIxvs/IOQQFMNf881h+5X+ywCh7rS6fDh0cIBx3nO0GaQkV6Mpf9mSLunZmv75JxmRkNbTq
y0g0T5Ai/vYQiJ3uBr5pdrBrXCkDKG2nS5XkwcOg21Zz7pBHEqI6QxwYsPnJgEExuZjraaR/tbD1
/qc/BtscLvicb9+2zeWuB2kOJCSGmit99H1mjKQjJ8ez2YkEbCifE/9Ya1qy5KHbsxjXh6rPtgf0
fpiwANUG+XBAsKVxYAEQMOk/XZeI9pzu29WKzmXL+VMm6kjhlsHEqlP75Dali7V8ydgRHClj2ldD
vXnOLo5P5Aor1jSQEHZcAiUdx8dlZ1KiKxfbz9enxyFqIkGQ7ZQ8VnKyhzVGqPnuYyk4U8ZGM4j3
aPE9swaNMH+1FBoz12H7lrUpJLr511q8t9KT0k59HMdNM/eC2r5B5/P4Pjj9mBVmI82rAdQhnyxk
7g1BgVu7SgZSHJVKsEIBas4UxfT5uPdcIl7oZwJ8FNWpCITq+zY2DYaRGuoQWIiZ6aCw3V1SQcB4
W2vbKmY4aGj20hkCtr6UBBWTr/kpaWpnvBCYMBe2fQMLWWne8TafYfAnhacDYptq0PHPWn6wKMV3
KOtkqqkH71UziBHAxWgq2yor66j1ietA1aBVLnEj7PHwSoZ5I7CSi31Bj9VxfQS2k8d4FIFY1MdQ
c0N2Cp3h3shrLUFITpdD3zzvgG1iEupwRHOAZucuAf6R0d19ixUW3PjW1RxhC/WZeTG4citekyGv
TU+95gcpFTNi3OYghfQcC0rbRZ7BleF0+/ro6oh+sc9YaJVLQhShxTZLpmfkwzjYRnUXd5bJgqXp
GiLHhjow79OJB+b1vv1OuQ1AZe+QHISgEikjgUA8AZ5UaTaklvJRefPAEBaWohQ6W0erSU+NB9qn
uZMAq435pEIfYNuYCHAC5nDgLxB5H8Y8knRn/v5G1/8W0W6G0m5gXo1V0SYc44Ou2DcmaN8IQTht
E7xv234aeakRmV5+xOrW4xySYqYxbjL7acDFTX0oPdpucI0v5i0of92a9AEzMP9B+TzKvsANFeEg
QYT+2/DL2SM4GS6f8rSXswQrZthhV7FsfIlzyAI29I+/gAdRnJE1YKKtC7mM9S8hhcikIvzf5JhR
6FvMPOuvYXzN/qVeWecowV/5TSKs4pm/++NYYaXz05sVvHlWjG+t+9hCs/MQs86TvOD769p/1PX8
OawmNINgnzfASt9bJl0n7XvsWK2iB7tXw0dqzoKR7W09UZVBaOFhemxMuYE7SxvI0oYZkOykdYZx
r64n9XhDnh46ORljBtpvlZ+uEYb2iaZULDUfR+pJXUI/V1XMNz0Bcr1RepKkuWXRoQa7OXjy+Zz7
UF8HNNiFS6q4vhafF12TQx13d1IZJD1q2CvwlESdO4OiWlJlJ6OWPpxFUBXGnwBieL+ekAhPiDgC
0TNJy/Q103epN+IvzMPAf6Jl842IU+RIqOQeAYz89xwasFwvMyjP570O1ogy2+bOve+OrSt277Sx
AT7GnNLyb6JjVDDYsIy+NNyQStJa4s2pj4oX6nSQEmeaej72Ohae1Xwn2VeDCtk8rwONSTRrANr/
WI7Z4lP6YgWS4MsZrEUo0DoT7j7j1vX7BQsB83bRbfPCnEpAs5gl0F58mEPl+9M4+YoLlFklbbCt
y0StYfNelY68aE2WZERrT1I7AWAyh8g6Y3tdPmA0bhSRA6knlPPhPQnQIQtL9ytQRNVYA5Xsy/bc
pkiJ3jdM9L/YKygzZP99VASRJ0zt9pU4ExcwsnIkpDDvskG8jWqtZ9Jr9QQPHCyVeEbCdBCkc8vs
UNf5hGm2BnGO6hMoEnbPEh26hmnuvAQuNlMnhWvch+8GYAEnvXmoNKiXLyT+F7NCBCxzRgAGcYww
IrlyoJb8SAKRYt026CCDmD69cHDiom/Pg3PAguURcjnZnUMGqKGl0rdpQR9B/pb8utISQ/UISYTM
+8kHbATMq8TtPS6k8XiHyRyxI5JwxFp/WwesMPhDgnphKxL7Kgnyrn8pWQWXhwIQwReN9sj94qRt
1JhpEaFRTrEPDeaw+iLtLJPYjCECNMTTPdkDw1AnaSmID90wjmBVPg+Z/f82Z7XA8jelAXFBtSDF
LAH0tCcn+mCqt//RWzRm0BGPcuAMnK3lA+na1PiLJLvjpUyuZx4CCtT9b0aN5ek8r/u/D1yQ7Ms6
XRoO3otTtp18dvmefg853aIE4YyQkjNoEhyhk11+8CRoPy3P1YzHTUel/J1AtUu8modB1Ni1QIq7
NgwbWAhgYao0mfb3oTRBpnmVSW/+9TRScMpSrICBXokV1kUNgxWWj7aQl8Iz0yVxsoeFf/eBa7k/
FMLUv0x7lR0djp8drRvJTRR/9GLTYpai6ID3SgOw42gf+FODJWUECKjW2iz+/vZe3Ky1KjQPf92k
v8OJnYq51ZXTbRVvMN5wfa1Sz7+2dcrfYPZoYiajQoI8BMtx73LmQ2P7bPbwXpFLiKM6us3+VCgO
TY9DF58trpt6G+tYU4UitX5lkGhCkr2+Dvrn1naaqVAroHKH67qpWatJFtyqQI6qKWI7LI0VA/Rh
OJBVuD45VGe6RzHmtBNzU2dn7wl2roayQQbn8KmEjiDPzKcwA4gHEX8FCKJ8KQ64PjMv27eKHC2p
PY4vW6eKeRxxcEUhSy6KuFqCcnmtVgSbaKjB0BVS0eBPLA00GkmPg1qGSVnu9NDh1PKELR60h+1v
LoQX1q+6Fuhx17xf7uZ5MCcFZWcK/9Z3/pEaL7ck9NlUW2dtIjhbzVVKT6l22XNkJ4vn8KARlv9d
7snXPw+uofQwhS+Ppg3a9I8w7Rlu5QPNsbDUJUcqhupuhqdPZ0avN7Yrocv2/M0XcTNeEapLcT0U
TNJ3aJI+LV+Y+u5jwISIT3L5wBMigJh5Kk+pYyM8zZfpYsF2ZCWXGfeKA5kVnfIav9VbbE3fzSjL
XgBqHegxaPo13YH9S5wJ3Uyx855JmT9GjYr2frdj9n0GSIpmuHeBo1zARYiEBWFVarDgzpL6nmtu
8IRs58XgmSWa9tHoNvbXyR42q9e8fxx4MkRCR4pu96DUN5QQpVmgrPWo708AoFqw3dEKe3lMEK0q
DFZIlv8M4cCjiCbVcVdIi1M91US8vNLK6otKYEfxggOoDphVXIlNQpCa5+z8s4drfyg0yOj6Jqn8
4mMXtJnSqn2j2JTWbnt4p3C4nlz1P7juI2z3QaghMy6jws3sgrdr9IJ2azhzZiU+l2FrFAV9B8EF
6efY0+IWfWoR4KlmkakQFLA7qpFT/mLWbO7+j5Yux1xRNfxzmQbdX0I3oAT4uncEezHo4JL+Lna4
F9IPSsQ1VvExZ9twArpDh8zdDucPliZmrzzKWkTWiReuiwlJTkWne6zUicMIGN7tXaSaY6GG5SzP
m0wwJKmcR0oy3bsf9JYdrQ8wFDsZcAtRpabE2/Q903C0CfPZjVZv+7ljBCqKW3a/i/SP/fiJCjSF
NXwWuT3KujrjI0fWaaa5pf2U+aHlnozD80Lg8nZ7W1hE9EubNHwjpyHsRqVcXTXa3DuuRZkKjlTO
Dr8o5Mo1nFfc6/gl4XlvewaJq6JXqWepGdXcxpR99kV49RpmfM2Z8jLPs6ER9xdK5vRq4Es60xFg
TGX9K91by0R95uhDwcwQmw5/w+FhkqA0MrUZLhwDsOpBMffitKa2dPQkx7XX/xvipBX5fbi5faOa
Vz8W4EZyC4zvFMFFxqmYdgz+CfLn0wVc7Ag0fSP25NqHtvhaE2GY1iehwqjjMmT7TIfUgT6/UxzS
MZtDGxKJ3rlk9rDZwY71LQRQwtrb1Z+KmVctI0MiTG87VZAMRHOGsQpN3EbH8k9jV3X/VU0lUhsr
W7i/5LghdQvpmUnMkn+d0WNZxeyBskx4lLapZTi5aQvwl0hI6KuZSGjZtdqhtHb0oIKLIPYvUxL/
SrIEn+YD4IsgDKmAhcITq3Z77kwCqd0Z7dstOfTxxRrMnjJZriIEH4nM3PeAc0MPb7sID4pWAAhE
unu0XPIViaRWnvAFImFVQg2yFbdwCCFwCTQ69rvQ/3lUlqU4QkKHuhy4z/SqrpFoNy3/2a3aS/fO
fH633stKSbkUR7aCGGb/7NcgkCeF3yp6xLzb1rYXqEOV1G4snqThq/lTBJc7nadRD0RVzTQ7I9L0
SE7uXn/8z1qLQr/pXXrYe5ZPegA18RqTCxYSPXfKnG5DK5wJlmHT3+WyblsHaSA8dnCi964kKxGf
3yi87AdRqtZQY+gYLjBH7TKcsa/AzgWYZwohm0r16y7CWen9q6ZXF6FXMvq458WbPidQl9/gtYiw
Psa2MMt8S3gL7ScQyhtNeWRCN4dzYG+xi+yrNRrYmtsIP6fhkiMbCpWfDmKosxruNB99vH7Kq1Pp
YJZFc1ALC5J+1fUndsGL25NStchYrakvKz6RwRQCd1CkwYDQGa9hKEulBies3NR4/QHaiFJBEBsW
owoX7xK8fnPgBd9xEAvgcz5LSzzpfb+96IOaU7mMLJMaTu3b0IpuwAo4ceiRO4xeuvt14xpebhvV
W4kawLMWeZOJFt5OlBo5l1c3/Hq959Gv+UUUNqLm2rc7TMvPrBJ7dlwcFFYoyQM7SJSxTCuKK68i
2n0wffPefqQYi4eX893D/Jw0hFR24IuO2/78tdpn1IEe6XJja7zW1oEVIoOS1j/P6AjkUvc7+hL8
+fzFYt2RxWCKu595C01sl/ziu5O/A77K2eoOqbZOOZ64GQP5FMkZWycmvlVM6np4imar7aHwsBbg
WkmU3ps3FemElCTNu+xArQoRkH7VJmKXfepRlhGWlOFlD25tGyeU3JoF2Q9e5AbanYWovTg9YMMB
nNJCEGIJ40CZZZcDZEHvkn4wxB69N06Xr+Z6Qt1L87MH89a1cBZQ2j5qV9fBXGTETh84CPdQazNE
jTLRJsRvz2DnBGgULqKbinE9YEy+k04MtbqlsLoNl+M7xK7KuH0e/ONxpu9GhC0zx+bl32WmUajm
404NspWCalQ8FkYNQpIt4XG+cp7UFsixgddK6syYNRrGH4tKINKrbux2O5zzY/cABRD4Vlwiyktj
SBYQM2A10GTK5FIv7JxBJP6avDptjagP8ED6KAr0Mof1K3ga7dqF0qm3f0cMFqowp2FGONmAca+z
ab8IZa+U1kJ8DOi3HOyIY9tHiOVNO4hAOz1iNpWNDfBu6j8+FcWcnenaVso8h55Y6Azr2WSAntkv
Re9bZ7v7QIbbbhAvnOzAaVWYusSq9t5UMfhZeNMvvl5AumWjPpRUz1FVVT23HkX9Qs6PKb47CGEN
uDEtZe0IoHp9NnNdMq2jf4syZQzIznEXFR8GEtS/0tg/AsuQGGzyltiQpCazFAPcyRzQ7ZFs9666
+xjWPgPngaQDv5F3Toeb5NaNXGIC5+8nn55Ta4sy9APFrI9eaMR4qIx3lDMQY5KY86mdGgEKG22N
KDzvIg8ip/gc0eE9EKxHewjqio3BwXX/WgpUuJfsGNA3bJBJXy8rsVjcW5tvOgQeNUqmqOJXyLFD
gAFY9+lulgLC3jTTT4Jc2Uwik5cT3ZJmegMIaNK/VncaWUa6iTSoNe0ZigIuENe8hCUNSSYt+Kip
yncazPpB4HN/GG43neC36zyIq/5J1EUy9x6R8vjMHHBkWP4dPNXcm+lXjuQ/rS7epxJAhwKqKl7I
W2ERqvQf7lz3t7vLqZsFJYr9ZBeZjUVWJlzFhn229/vqsyqGzh3bryNXWjw+UgnsuHIXgb+Zxx1d
4fWMrEz1aEreSqXI7Yzkb4P/OgxLHvZmkCNzB9c2GQLwhHIa8lyGTFEscH3vtpty/Nr6nYqbndmv
bXcDZzq1QjvbVeUyG8KEVGFYl5QAuW+8yVNfaAcFGqsaGQU1PBQU82dbpCZUtrdmczsxe2/dt+ka
/YOtqTplkqDkg4e5StgB3w0OXun2ln2tu+HwxVMm70co343styR4ISxS63DvYS06NgnzaspynSSk
N4oTo4oF0Fcx+WCRwCrlJKfmloqnRQb7t3Tw88zik5Cmr7op/XAQ7HFOiG+K0DSf58Uc07lCcfzk
VSTx+vTabURNJdoPGsjRdHnlLjKDvwtmYvl+ZygCtVe8NAeMmsZAAD2aeDr+gIbkAnLKIiYOcTAf
rqmFgmlSracMQr9wXehuLucDoz9CU9wdaol5FVH1OPTtWu2PCue5pLb1ysh/55Vgo9joRDWTX/Zl
n+4jxUHknHvqT4/aZ/0mAojomy+bk1mXRrNEgAJn9sMelfHIKgamrRcS1AJm2WIdTJtkO8WijpsG
ldfXpPYx2MLZSpBQwt2Sl0/ZCEItU8Qyw+brx4k6MFG1nMyUtIPCQF4ThwkHw8AWzZ/aIMtf7BDk
vz1MOdXwz0RxfAAQce7YOwqUlrRYHC7Ti+9ayrVvUm3UJp3z+X719A7d/iDOh7CB+2fwZPDsXDwc
JLCKGx8TpmOGm9aXZXdlY17hdUgKH1f7MJ8VTR7YP2MNYR7zSOCMmv+AJMSqz8Vg6H1jedvtpWUl
TCF8jma5PzoHHaSwEBLmLUr0eNRa/JlXO5E3z8LQXLgvDKiJfekdHGZruwyFO0KmYIz3OVsn+752
aRPXFcwNG+gnQZ+lb1o3kEqnWfMHQgl85Ziu+mxW4pa5jtFeN8LlHDrxALF1rYR3ooKb27aKkv6t
wTmjFgcRn7OrR6OnwJ4whi2bKcUnu9rcDUoOZXgSvRjWlUcaYchULwX8CfAW97QBOelNM0lmpFF2
Pl8RRKFUm6vIGmXT4M2OyfB3Zyl1P4hqRlsC8uEOIhV3ntOScDTpQ5Pa3Ap97eKkoDkJ8uv2qXHA
OgfbPJKP7NLI+OWkzHdyIRTo8UvFkNGPO3RCEvFoAX0cMPyy2p9Kq08Ty/jm+CfzbIu1KUFBpd1f
x0qOPlRtF+04cwVNbf2CIQynS8eCPgkBNmSwZqFin27ERPj+jlojsVnhkBx+fSBYo2LV/GafaItD
6wd8vJvWu9WIFxDryxXPRR6q/I2oLKj1AHQHvDI7tPVK6gCF3NIZ/3krCrYSKNBe2Ldsax2szhEh
jkr0p2C6/+ljbOslT1/GrG39+1WY5ShYE8ucOjOLtUmKknEZjSIYhJan6uH1lz5/JmAuSx+6+SqS
2Tjdyvi8EAXXOSllks2tYumOxH6FAEBna5s3VOFiJX16RW+LZpJgm6AUhzOd3otynZPU+cwVGlCY
cttA+c3SPlYE6zDYLDfBREAjaYCRwSyRma7grzyHvDdD0Ruw0tyDE2X2Wn29b3g4PQM8FgHOvBKd
tfKzpPsXZTa5gEGKb9VzmRe/RdZ9STYk503+fcTTqcU3U5gWUap9yOtBF2j1RnN3MRVqM5O5iIyh
Qm+6+gjun0He2iog0RCkcLP4mfPwM7WWrGmz15a1zll1GbQ+0J+tmly+Vpv7ZEzNV7huhhPwP667
xVx3I3dJzoW8QEXg/+nlVAy6IqM4Ty6tTCKNiF1RoJMr116mjwZIADtEYY/xedmQP8kcpfbvH/Zx
eg+qN3SWZUMFumnEenp5+G3J9hruVU/vS/H+JBup/7YZHHij2d/qP9jbE77yy/Nhf+anI0eBRbHA
dOfmOT16aTfbUK37oYv0I2R4gxb5vRmR23AyER/9ttfCFbQK89WYnfMNcGqnZji1Uv/41aI34gd3
VbR+44JiiDt8YcfH9BqY+HqcRHJ3EzxsRKoDg1wF7DN/WbSwfVO7RyjjK5JlCymQDraC6VbjgfkX
VP+uT7ckGTCzqW/B5mZ+1xc6a+6wvRjnBqvwvle8UbxPmedUCUbVH+vNGWJezP03SKXIUVtE8w2f
uow9DMnZQQj/KNh0Hhe59k/pNjwzKIh/p9Plo3PJVZHzT5KFBoPwJmvSBK/A9NiEhMx4MB+LAWjN
0/heQlVBsx2NDE14s7fwGHv2hFEFxqNCP0RqxEKaVu9EcflOrTMhzn/G3Snuq5lawFJ/oB1aANUT
wIUupAuaGuFQDCVYLqph5KZhv2Q7dIyHBzWs6uAJ61o7j3ixoxCHzytL9ue8dhemcVVX2G5gxoub
/LSb/0xcsnkJQpV1QEByYdF19le6Mig1Gg03ucH4St0iDfEL/Q4PwEbAuywt4cQ9CSxHJEUHnj/y
AtYDWbi55R+DY1L6kYudYgYYznDEVc1n+xDph2QufyD+1M1LI6kOKNBg1eWi2fWfk7MO73aqqv+d
FPKExWVrTLGmiySbT0Xk+Nw+R9q9ZbCgSysH2Wjc/oDn2fTNhGQpv05zj/5FQpVISa8+P1sFrqst
FoR8D4k5Bt4aG9fe2amWnVzze2v9+KRJZFiN7wPKcNTcAERtxDyBB+o+AjC+WRj3KSqJc2up9smL
wauMEkrVs3Uh6amH0Zac2nyz5auYqIAoLvOJ9d5OIeOxaFpf7X1ixy/CK+ncPOEgpjj9JZX7UOEg
hECTDd+iIcw6kEhb2+haEr9w8iQSFEKB3yXMxvsCXqPz8DkbJ4xo5nqQeoQURPqSQDYfBWpq2w1g
HsX3/L+sI9tFtW633ApQ/iU4dFNGPtdxJ8b2qdD3NwODE/sUbtX9U26GEWIsfKIKlGBPBJAKLwfV
2M679jg56g7cFb22x1+mN5EBQV3ObINvOfD4yVkTDQJU3SUUMyANpbFjvIaZiksQKH7MuFzNo2FY
0iXWJGiOsDwBIn+4Zl7xvOq5IGqgh6Anr73k2rzDvdM4YAmkJe/+FpAhDdKKMrX5pjwnnxbI3fF8
7//4fKBVh0qbVZUj9cI8FSVSnwtpL46wIoewXTrMKLYQfXrQqp/Kvmo1Naz2B9/RlYicyE5qdLuH
QvZccxHv9Mq2dpcJ6OXjfIIExVMZrmjO0uq6VvdYs44VRe0utcot1zGVarAC3BvW833jdMDahD97
T4fuzJ2bttxl+J9BHCgUCPgCD/r0+UtPj4+Tem/itL97Q76n666jc8v6+jJdx1vhKxbNCupiai9c
6CHV69v8VOMBhf6xBzlSkmk5U/hXhK7/dmbNMzA3ty5MZ5nADkyUfeJgyEQyqwzly5cghxR6eZqu
x1d9jCRxNv2Y+KElRV+szSulXqHJAYPlZT2/DZSdWdOr2n5bnspWXLqDJ1XcaJDR8ggBmDQBSDA+
6d7V1WuKxiWv3dxam7x+LpQ5bLtUotlAUH4mhpnh9lgs1ve1fyevD/aLRZO8dYL+2sa7hyll0tI+
/46gHQH1kKXsjtARxapZE2cp4tfAmZuTycd1aZ99prwzhEvjjm5jcOCb9AkfzWC1dnrcUfDjgKKu
Blv84fUotD2MrIae/zdWd6lJDfqEAmXu8YESsSs+6Gg9TBzva0SXXhj+vTNnV6jd4P4hxQeY5vkF
aCVGTMO7jVxC0HTdQYZHhgJ5aYfWKlIQBRCt76YBMQGSqEU6UGEzpGzFKzww8grdmde1229BRHob
uGNJ3AYk7DAk+wtshNBpXfeKQiwbPHsxMBaY9IoWrhl+UnBtgfL3WUiRoz5FRFYOoyJpVnYk9YwD
1EyfXBZBfZo1e1V/sPgjJc7omJF8nxvgbINoPFhWA27gcUbb9qEeeyKS2s8Fq3PL66W3+bDeJjEk
LlHSgg+V+qAk+WaMpKRi/g5lk8fHDvv7kOEKx8Zp5yHwW3TE0Be2t6BfHNQ5VFukMP3OPkpx3ZEv
2Hk32k1QUkp3ICVNl7LRr/TCw4SF4yWsWxXmxB8rK8Azdu6a3K/xO6wCLV08eJFYjCLNrVyTKZ+C
g5IMnoxCTNXeac9Gpn7KWj7Hli8zfqCY/5kizNSlpulGd9WdOr+h8x5ebZdVdMeRpL+pDv1hv1u0
zCm5dYLqX71RW9UlSZXRiffpFf4cRRyHhEE9iVzqO3g6ioecCMN86xp7OuJfqiyLuGxNbDhZu5BR
xFxWOlZICL12rTHiY5CSLm5otlIHUjZSfiLBtlm702h13+HtB+30qZvKpp8Vu2SpojB2jd+ys0mz
7hD7acRB3SQfigGjXF+Dk6yd59koLDlJetrM/YPQtkK1LCt4CKM48CLaeU0rb/NksJuI+uc6Kq5A
k923vtAzXCTkAuw0qG4n8AJcnlr17G9JcczvtId2SGGWS8UgociSh8oe0L0hU7ouEyXmKPRnxRhm
X/yNhF4r17YVTQqL3JvjBCZmmPuYNU7sQMLsJkkthda46583brLYscgnlKkGQjDbQAF0aaIm5n8s
82+b8s1TAWfph2gMBE+TFyzCpzs8A+oTD5kpopEVx/Gp4Db/OAvrPqgOvVCkwssfyruqVKo/3GwL
0MtaAaDgQRzhBYCORrsGuYqY4RuT7kBYtQtXxRPTktvG0Ewa38p50sA7NNVRvTy0IJJ+p62x6kVx
h4H9b0KLyjrb/D7kVDv+jYhgnccJxc9AtLp3Yh/E5CBx4OLnKSOxlvt1R90QHbuvzCn7apQLnWEl
eyJzeGM51sZJCD+8GXnK2p2b6t5ehWcq+SqT2UZQs1FBh8fY52QMUJeKwLTIJDrE1wbElBER4ddl
XpD3GbY+qLgkk4/x4MB4WmeERrV51M/8tg4VKj2ypPgjHTvXFTdwnYCgEW5ySofdD1RYlmXmp2Tw
EPT634kJHAs4ZgBGJHoceW5RIAX2GQ5WoJOmPWapa0KzkcbXt0yGDZiDpVmzaIer3dcztZF2ZyfU
WJyTZ99fruHgOwflRe/GrLzfDMN4q3VBP4WcjnpwO1LSUW6+wo/XVWy6dX8JvwV+5+/6zCCy6iw5
fULexoQz3G//YyrGqb7U5+Mhh2E7z+Zcvw9PPOA48NouJ+O36Va7B2QJWQSTHp1UmQD5oNrZOspt
S70yLlGfOOLgDteBWi0YovXoML2kMbHM7i7vRPa9vkrKr38wLJTIDyybWSxFImsAlhzfz007eg+g
D4QHdswSXI95myJTTzLKaSY5WAof4GAfexizsCFZBo4EJ94T0YL59Wi2crfMBl71unXxT5z1Zy8A
nopjmxvHhWXsOeLpBGLO4CO62yGoiu0LiLoao6mkykqEhuBlpPKDpjDHcAFS9grXJP7S7CwCUkc9
PJ3VtwzbZub12kXHdShpu0a4eiu4CdX6r2UWJ5M0JV5vKSvBwl0uTQMNN+UrBdES0IGbU/JgNui2
zeYJJdqXcBL0trpNPm7B81XiAYPQ60auEHZlAxQ4M7hxj5pT5fLhKZdzd5ul3mjMD7f0/6Ng4eqF
7WxYWvkBk4aBvxiM20cFAxl45YixSOhrkOldKWFq9qO05GFkF9m6MRCZhiY/ozmQtIWDUw17e6Na
GZ9hjyEyq+GOPvL4M2px7F/FlvnejJ1raLIzm01IQ2dICnB37Y2Ur77iZpwR0/ENhW/jWTCl9V6d
IfyIgaTAs0wiuchjMGNVQw4kttqscU7+G/kj7xfaL3HSci1YNQ2Q8E4lCoPulyVUUN3NwCKW7h5P
5l8vDivQcyBQyoR8G4uE3GGIh07iePyWqt/MTfDRvdqmW347LiS+uxU5PUkb2uJVj0kzBn8mO+0r
Zj6vN+ATsdJ3B6Nx+8wSbN2rfV4XgdzmsN9A+muMilF2K+a5oLYIWMngYEs5PcMchDfILGk/aZt9
GrNba7H2eQrtLDgew0ofZiUbLRyxwTruBY3rG8R84zAY4D5+KnOK/PZKWpyBVryvveXQU2qX/3or
Nv8ZmNIA0GXvVV0cn9r0NyD1Hr47CxJxQ/DRa+oNKml0aof6xeYxJzxeUs21Wl4/S6MnrDR8LHDw
XX3CJNJHHWpk/6C74b/CE8SfA2OGZf7kHPgODLd4wOosj8B1B72zvX71IWaiNqxUA2C+5Z3uNb+o
UJWeAWZA2hVUsCFhOnpRqsZbKGm/treROBPBGMI4sldNDXsiRsRtD7UXV4Q1vtN2VDtjtGPyoFBX
eMuQG+jLxBD6AuhWsfBZCvfKMclPZ6j899doWKENYdLofXOZQQ6IhF+KaIpzU75fzvVKsoVajstp
P8jgslBP3XVB2lLz2KmB+EerRwmxJhAgWWkjv6tb1Bec5iOZmfUtmHeSjuqlw18kQSh+/pOrE+vM
ehle4T5NOQu6rEbYifdqpkU6liRwxITL925s8AiEj5+yPDwb9efOFr5K+/EZDSUdbYDKOW2c3g7D
Kwd4yhPO8vcRtSicHijaXdYmx0cg84LFnbg/DfMOb4Bk0E4jfoEvKdsmxLq3+uS+97GvEHWn/3jv
WCdds3l1vFoIgCG8a8RlLxfl0WVByJXaxPw9M1Va3mAS8Ptz9M+SfUQse59wmW2ImzFT7KkYdtRy
1CciJ7g15M+6SXhYyH8m2y7cylnG5FANzFThzuBsbGzQMKOUnAwH8pFZoQE2bvCiD7zLF5c+MoNf
jSg4oGnZfra4h3oXoY9RTkwACGbZ2fl1WblPN1+4Rti55xO6rgIeXyc04+6jO2n6vWr+VSWVw95Q
4/orP6OtQ7QuwCabbmsyIwevU9UnQVttgJpd/XTUKUKpceHEZoVPhSsjyRWsavg+mRjBP6mIRKbt
M1jWPwVsMx4jRFioLHZooDWLVGiLy3UXOKjpiEKS9ImYeMwwh9NR3828X0j7YnnLcvsv4WuikZc5
LgnppZAndAzH4oEh6riYzKT7j3vK5G0bF21v8HGaQwPdEgbZpSUlkiwM4HHyawm7QUnO9efuAkhM
0sNOTa5ysqUaPLSC9T6MPhHrczcIANvD1+SoD/0ucNGpOBX3hK/0f7HdruGZ8b41wsrd+sAG13uG
7Om1B0vnMHEZUzdhoeiY0CmlqGl/LNCbNmnFNMFDxdcANn9ZsNF5p8s15VuoZE7D4vNemT+b11zR
HLWc7jKMwvrHdjiE73fs5xHK25aG7NprX9ttobUhSbnK4edXbXLjk9UUOk6AttlL31TVd+9H3Oxd
adtNphB6WKF3FFMHV3uk3ilyiMMkTDP02WHflhk20MtoUMX/f4XHyUWfE7UcRMVV2yUd1/tjjMDX
Qu04abeDzehv87qlvlfu6f/E961dgjyy43M2FAVhyi8hI2oFlEr3hDjilgUKUJSSJlw1xMsERZKq
bmX1K4JNFC12hnx9jtBU3d1JoIozARIhwbT+u0owyy1wIBzPApFP6JgVXJjMGLTME7R+GXLF2PWV
4ct3uzZfkD63yn5/WA724mrUxA5e5Yo9S32mfd78EI4fgq+LU2P3QPHV9rP7M8oivW+sWbMD2NaK
0y+kZhw5hE4ypyfVAoemRrZPgxa/MEO5iUjMK8+ods3ibwx9S5b8erIlCThp04MD6ltBXv9zYk+7
wdpUuX33lZdnyFXkAixR5/XmTlKtnDnSRnSUDGoqLA8zBFyGNa37sKGf4MHiq1bT87zzWo/SD9Wx
1q2SwdAULMjlEShrtAKd92G7vVF3hYcZ35486tlIZDM41auuRNtm2qpHNmoNMu8KZlior8s2mCJo
217Yf3en47o9za/ph9/hB8tw3fAoXRNaXQE7PhSq5w4kxuuW88yCWPCxx9mvNg3f1h28yzYDkblG
IxOSP7GErlaUg1prbCOsffBl6fKURtyec3y9CzNlMFMPd6xyS4iTB1yImLVoqvvdQdB20UIO9Ggv
Cvwl2lMHdQtSP5csRmc2bB5PnF2m92d3//d6pcbPbUw/006RiX5+45dKrhPYrNfHw/XYpRoaWI2s
CR5VwoASPWTEepjPVDSwMXLeFSoGU7hssHQfJR82NlDCOnrKoJrjpNFmcwPjtgsDDHyStq0RJXyO
4ZTgjA57cOvDtZpQoV+si8dmqtvDWpix87gOPjahsJ9I3xkOb3Pzz/aqE63wDAKvTTTckgvNZKie
qc8AV0Wq7DZkX1qkbV4tORkiUkaXbYLtWK6+r5iwP7yxKAzl19pVnJMI6toeOAkvJ9+XC0kjTwUK
D9le5WRSf28MIdWFDjfzYn/r1Z5UCnG8Veu8piewfQZ2Gf2DowRXydT32vdN3DTdrpIsKw0y41Or
3EV9CDi5Lm92BdYqPzOX/lgS7sd/0I3xOgiNrQn2YOf6yycjmo6uulZlXTSoKPw6ku8A4ilmFGJj
DoH5XuB5TKcPcs7L86vN7mVoh74ihowLO3ntLUeybQPZWveYytKE57MzU7weq//3kFXJCEP48TXz
75odESVAm9NCD7C8RG5zvCCg4qtdkp2qGBCWhw2IZGNFYOXuQfRyZN90gJNXu9UGGueu0ug4+clT
hor6ykxcOTOI/F71VS9iJEKJYWus99saXfraLdonNpjW397omZfbWowxkL3LUio7YVr+aZzV466H
BFHtbjNhqb4FCXAjDeFFRGCCbWUTsH3hFCcieS0ukKhiq//9L0unYW3GXwOLp3IBc9d0G+OU2j0b
0XeKPAEeKNQPZyY/mrF1JirGO+0qgphthTXIP1IMZP/KSwCtzfeOJYHHEUMUdUsj1iXEK2NLDYQB
KjfKG+wuxTWbG+2VTX1wusFTJ/lz+t7dZxn4lYi0LCAvHcwgcaKaI+JphCqHoxtzrwfAH5aOvk6D
yfr9gjLTqWPSDNSfMBtfbOvx+0HP0CFMsxi1GY21hdmzDDCW/q7MGlbClAjn/ffb9cCw5l5FBGo0
VX4v2vZ3Q0rSeEp3/Vq8R7LjZ+CZYQ3jGr395CY3v9hPtzCKJW5jj0gOJ0kko1AS2zsO3fz6mEXm
iGVcMeBqwXMQJsflLJJHCRGXSJSrYJyheWUXgy8pzPV0gssDkhK2GzRzaW8kvOba4H72J+4pORIX
q4P2wXXMSbz9uJKBifWZ+ZXoK1R2uBWXxH+qEq/rsGE7IwmfQi18A8XRP1sZ8VYw5IodDJilQIsG
zLHo+zikmr11jNMHnW4AANvVi97FIrXh10rWAPf4PXh0bU8SULU2vWLDZYI7PLTFDctHlfM3gNwD
6uYVo2W7uLFe23+/5zH3y0U25sDwbt8Wv/nN3SUD7rW5bmMbUPFFOmvc73lKQO5xI7W7J0EO1CVl
Ha8Zci0/so6F9ljqv0qqbCWz5smV2eku2zH6L/JWXxTMHoZMsJQtxI/FOoOjjqZXClYgJGiCRxHZ
V0En+FzPtRmgVV514bt1AUV5LzfR1S4QsueE0hOaP6yRy+zzNY1Mmuxa4PwxW47lVDtLL0WhBxGA
giqIrDG2mqpXJhyDw+61izQMesimlXvMPzYy5cfnBLr7mItD6GvKHsQBSpHuBndX+X1R4JkPUU24
nj0xLLPKBQ9meUzax2gDcWgAjk4uDzJuFfjihcUtN81fXYQeKJRuqFi2jtvATiHg4szBu9cDWTNp
dPCVT+Zirx8j8PAFl7ljHR48bLiPxRqZVjyuD8IfcrlPN9E6y1mngYkiK/8XACTUDj4GRgZSy7mQ
5Zpjcr0TfzwZf7iRymtBKhyspa6XIkEzpOsm7JtIhN/83ZX5rl1zgi0oeoVgtGTgdKuJmPKccRF4
N15Kv/UR0lVrF8hK13KSvItlvxP++Dg9hKG9Hh1uEJhrApGLyaR9NXsBrZfpT2QlCrmK3qSidzpk
f7eVz4C5WxcxA92h+/mwH3P2uZV1cOJaAvDB/S8I/pvjfrPCn1TUvw4vB6QLrXmvumXLgf7vpemC
65wINbai6KRGgRJSBVVuqTkiRWeTxS3m713OdUY7lge+WKQijFHJ4pHfQuyVtdCQ0hvV2PRul2QV
/NrvtXCKlL8vhIEjeRwm7Kiju8xGK7+GjA/+YisbLvf/sIwtFEj0+hlnUFjoAGxmjaME0e3KyRdt
blwVV3OrLxzDaNabJBHnekifY7I90HD5H3ROYxbLtS2Tk+NoZ/CSESHZ8+j1XWMLyWZcxq0cMYhO
NCpDdiyCBzPbMIwDJzcEYJJ78gAj+kjaSaFp5Zk6yMFiQMF3JZ2RWTlShR/nyDTVlNa68pIPNkFO
H4zdyGNat+ZnN/LMfsTM4t4twVidUoqdQHYEZVZep5OYyqhwowRecnka0xDrvRlYrhDAKFzNbjIu
G48dvoD6s2VwJDz6/Ali08ktwz10rRy8AsUMN3t5CQm/LSjgS0yR99xuss1Qal06fTRvs/7vXRx/
T7GYJnkcMuXZvyAjW5oneBM1rkbWVBfuubk8IFC0q79DX6uakRq8ko18VgPvIctnWdHzs9kHLxnp
yOJ/Cyi1n+6phhzM1gg/QJ8MceNAqHrGd24GLmaoK3uxWrLAJD/S0S7aaC01BlzzxIMJLOY0ixvn
lI/pCeJ8UtY3+bBgoD6FJRox9g04USUKxblXEjkQ5A5BPI43fA0RmjzBCBHXaqxZpcI9k5pt1db1
Crn5cxdZLcYrIi6i4OvST7+ztqMSVoF65RDZ2+Tpo7aUgGeMLXwvpx1lRaX/ffdrWK/7PPF7+ZKz
+v5VULjk5QeErqSmsx9cfP6fNBS8FXR2XX4ZkshkevUvTYXGGsmzHKzzSieCAp3YEhpzBnifP3xs
tUU6ZQbxfIZ4n3Zqdkk/njdv24qnyNtygIeTS/Rj2/80yZnwYIBkGO2hJAeg4EHwJj8wBEo9MsfH
jmsdbpN4AI1146htTvfdlLflQQqq7zGFoYVprD7DxEUJmtySSTEfS67D1gGhSM+W3aMrCNod3lus
Tycs+tKnDCDyDPozBOIPsRRnleZUhihFkm/DUabKsTfFRv66YRLUqdqHW8DOPgVQxHgCrnCRMHUn
Pri3FcMBZuchvkaa5QRBut5CHP4LcyOEwgzTh3DNrZYFO0AeekancCYEponfjF2bWdymrOo6VarX
FEAdlib+C9iEeRQkJUxZRVPEczYS6Fgalyt7CfVR/xOO1Xb6+kG3lHZZL/etRfDY6RpRBd2H2B5S
uOeWjef20p2z6cv6RtwfUmUnULRYNVu/gCgBZoKanI6ZLDK2CCzgC9M+7/kmcPTN7C5Lpq3+3zr6
Qx4I61Fjwyhpw45smrC+K6uRyx/nRI4wmzYB82Epwavo/5KBWee2JZ0AaTdgLblYosWySl6aCSCT
UEFmJRWe3yEdINK3s/03Fe4O/fH3qQIFe+0ZXUQjvKKT7cxgibpEENVkqnUjMiFu+2CVGeztla3U
aptQIpZSghDOVmssA7p9vTeDO0S3t/YFS9mwJVBHi/0WCuCSGiw5rq519ihkqoOo/pSIpMnsA6Dx
YuhPHcqI2+lzrrjdwPU/7B97PqlW2IgYtx2ajvDNvIpPB2K6hdniwCLbBZ5UwBa5gUmXFJwCZJT+
gP3/bzALN6N0iXdKFB6hFcv0QTOntO4v+o7Fb/CLzYKoxHLHg6xSYIU1m1tw2EhaC8TpOGR1hwWB
GXPlYyeEVOkG8AUjkvBcZywomIoHWC+9kVpEo6wUQC4UxdAIzK5PUjZNJ/EWWCJcr5DEB5VltJ5x
tFz/rZKMbyiqJUTIJ6IHHz0s+/3Thx3cmwLQHku7r4m0zqt6kRkFnoorw0imgotNX5+Lu/NysXC2
QxABJCkCUgSBzuyC7bmLprToKLYsSvtyyQ1li1AT8CTgxiDSrWKA0SDR1jWHHyZ0QkqtzIYlB4ni
XYXSE+bTDGsTcw/APDyYy/XIXPwjr4lxkp+Svi1vmSW0+NHKNkbZuJzdc8rjDOygKen+pTuCIQec
C6yGalwkJdGxYdJ2Bs8zIxxErbGjuKh2kaS0kOJf1zoDgDNvFEIm9aWcl+FDnWdjkD/pwTHkmeOD
xso2Hz+3/OJfovAx9sf5mUpFuDIQ9X+1EJK1gMk3P5FLPsgY2TgXKvVKSsKfQfWNFWY18tvWKGbT
orWPI4H5/AEaLweAgq2rIEw7645kxLMeAvnHePruVwWzox11szhmf5u4WZFllCEUBkTZ9VbnToNt
o2jCuZfNULTKwEBvhMr+YNlssd5yrLFf3BqJVpQdbcpcqAGhlANB4qGb2fqq+J2dQ+8uCWUcz55n
pEvDVCxiALheDJptWygbxD+xcR3TK5TEwqSva+JORzxTUio/u6YnYTwwSiin75frclQd8HnDBiDz
AnX5Ys7uWAnTlm5kN6KeyiATryx4fC6lmonk6SoTnbuJgx0o49bB4LFqrOwbo1jqMqDBpQCdUu/W
g+4b+hHz+eEvekni1af4u3bsevjtfXHJJjHqxlE1kQE/t9HFmoyuJR6rzNUVDCbyRJgSCan2jqpq
5j+1rWaxNutG9bym3Yfed/B3HiIWeC8YwknCTUR3bCaAlEGHr6EmMp1tA5c8aIZ87H1JJJDPQisK
cAmgggwu0BxXie0PMnXsao2ZYbHSCDGqGmxbNr25jsKGZTRa4hefN6ynUoJAeusKQhEbck803M3r
HEo80jRCj1xcK5OF6mK6+9ax40LwhySWB9MOMxrLQEXmPxRRGGs5fc1Xtf8PcWFOIHM4ndcPbXFq
bKT/BgJQTvrcE11YB2d1EeBfRAA3cOVpabJjICMQjt4k+Ri8KTg2H6+aqdSTqK4jnF1Ln6Hi6nEf
aCISZAKuFBjlduW7yuK7m0MdP+uMh+l2Np5fCJzwjXfag/iNu997lXYXbOqM1H36uUem7KMN73GN
6F991XvSFtpyWsYHZ++8PnnN59spjpjLlWg1r2uvD8z4KzUEkglD5nJ2Ku5LyqvvyIb0cLA6npbK
cabHpVJ6DwvLeNz72j6ZDFlSzKd2Tyb1Vg2Nl3CeCfdtVZszDGVqpCDWtW7kEaLYBqsaRt5sWZJe
yQ/oYWpgPjKMQnHBXBeuTVBHJ71hQKBgnRjAPYjBEtZPR1X5cjNNWogVEu2VJFV0KZSQ6S3frM37
i19S7zB/szwj4GSr19wb9EcSvIEYrIc/kBGqsXDKUHfDrik1uXwP1nYJaH/omyhRiDlWmWAlcfQi
MMVL6EcBfYZ9JMfSgDodnJGElBgPWxnFXGfs026H+9VBAPA5jFFcCK435OLRe6WRAOA0aJWE1weo
lLyGoPXpodgkDjtMYZsNztlQrSA8yiEsp4OxU47MQIx7Of3OEXD0aIv4NKC4lBYuoFhm4D8xTCs8
l7xY7liRvft/UK92CoLOrc1Ddb0xdAYA+C/hCG6CJnpAOZBmjFTTHiZSr5OiLamjKIKxf+6J5ypz
aN7Xrr9xJ6cywHsoPPaq7Cv3OaB24PCiVNRxpOLTiOohoHxL3P6iLLZ+0rvkLQNKyHv1T/4bhunQ
Koki/65kP3vryzbBSMVnzGPGTrT1ce0lUf3IvdiSaQfh5BKv73Ln3VQ6iKo4NXzq7TAGZcuw4owj
Yu98tlvfzS5Pmx/9sQ3U1OeNyA+KPZTeGn35PIeRl1+imgdNvHhupRPagMDrXqDMKX7sp4kYgw0H
ooAFgRZWE5HtpjpDr38wrKjYjl5Kg8xiPkWrPt70yeQ1Aca3H0cMs98i3UFfNV7fK9ahuNodB4nF
Sxn6FxGdwhYbp63AsGAbM8zHxPIEIthUq8mm7htTLqWFUGJhJFno4IpzOnAUmIsaoQ1d56VQKsD/
Jpe1uNOaEFEkfZv/c2NSftgjHD2xmNuYV+a7mzS9ZyVALpb0+C54u15qWPsM3bhnE3FgnbZ/yOeD
Qwx/R5Sl3Sh+1vknicbZoxsA/xQ1+DjSpuwlIF8megQ72ZzkOGmWqN1sc2sN6J0lW1ERqGeZ0uKN
TYs7D7bd6abSNmno7tCcxBFYoFeyMYRaDFhMA0OkCRFV0ZOj96GglrY5w9IIliTQjiLtxpt97n6E
OF44WsW/HFO7iBqEz8gXdV6VS1LKmGzm0bcA7NDmHZfNrgcSpb2R/NYULfBxeJFUepRtrqGUeoMH
TEC0/JTae6jOo9z4v8zUjLZi7Ypg1724/nyZn2fxCFTqb8WCpTQrN8hzqoT0fcVdkOnz7xsUD0bH
c+jEVH3y0BDaSAO7QBPvWLPUV3hmfjO7FBczxay6BCQx2kYJs/GOhXjcVgZhlbC1XpvVGDcbG+pa
PFmeR20wIJ/1XQDQGwVuPuHLhEWdsWs5Go003bLurAC6OclCsgUxjY1xkwf7cGlfIk+WlkOlsS3P
tHGOJZ+yi2rxl+NPPQGL4Y0ETKTE/l8iQAtOF1MMyDN0z3ztJ6Zu15kYaW1A1gL+2mMVtWSsn9Kp
MveyaC0HBa0JwzhAOjgmBn8ia0Xf+/tYOejfkjjPzGhz/89TWBdCleIAWZ5ujPrYOw3UNoPPkxV0
2oEWFcWRGlAaEONywUFDGIOxHoeYZnfcoD0PKfQEZRe3R48dbUAij/DSszAZ0P8noLVJcK9uEAUh
bBirwPLkweRHkDsf0vVHmCQzN0osXGMaAeJh8AneEzdPGvtFb2Q5JLlotQIIxCk7MArWDKfmXIZG
+WObwuyIcbRC5p0IgYkU0cKGdGsmwJMTS1kUrWOIRifXGT2zLTs6WrEr2JLs6w2kNEpptQNpX62a
EOvxZRSh+vvexoFIbP4AQXyQffK0ng6RoADrB9fRw6THHls/fyPw1SZJQtLwO+orLC03yzHOq96b
i1A0jGmE/hGcLKku+L6FBYlaBV3y5zJnjH5Q8LgiSof2goY5UaVtIKR9nB6/RKIat6Q1Qs1EP1Gd
dGsQTBfNIzLfJlEvbBVY77CVtJvfqFP8sIt9AhBgcyXsFllZ6UjTh1u5Q6mjZxiJIJXg+jyqFCdk
GxFzUhGKJD+37jwlWVdzqdM4SiEgizssOuEA3hlCJbmt0JuVtg/T9Ic+Gctt225v21bbSTxYaR+Y
2Vo/FFiFJExMgEF06cAcPr+1PLc30GrldvMiZCNWebLSbdVjz7Rk0w4eAU7iCtLs05RDiQthnxv7
SrCXOG7Hbc7/GMROSirf5sMZcvxn9u2/b0NWvM3CElnx8cBCZAE8vPS/yu76mT2cf55gVQpD6o1j
7ldRuUJddeezs6T6g9kzJ3AkrzrwhiRVdSFZqWZtbltZ/PwFekK9hB5FxIMR0G3IA3fyCL4rG6y6
KwpPv8guuO6yQh1d9799/9oCqYe8tqXt6Wk8CdQr2I7GRESw/6Gzc/emRW2XfE4/ZJFSZs4BU8b8
JqwncUvYAcHvSDlGXxdnEqNznz0d9Eh2K6wYzocWP30OP1xEIGfBUNAEwjJht883J0hZc+fJCacy
mTM+WcTbm+3bWkxz5Re0njWcxB07aWp6taS5WT7ktnkFIixGsR6e2XuFmrsAPVsdYpPdWoi48lhG
tIitMVF2uHXgIMo246cKWc9Xu4zwCFONSI+sLER66JX0m8AfHW696QP2ahRSwHCJUgxvPc5c8GQe
tt7hkvzi+q7LrbALWSoRqFu4UeEIr6ps9WnmrkGjvNH4NdupqSDD3zPuJWJW+vqeJm3KS0APY2Uw
ROIpuCecghHp16MAEykMlvi7gKFsR0eE14kvPOQJ1Tm5nZWUAwkpfFRk6puaDtOaMNoNJtbNSPax
n/i5E3Msm9+6LJPPUv9P9R1meGdEqBx0ptlkC3njkzxVd3uqw5NW/PAJRL6UamUopJvXiouGmhv5
rNMBlvI5t35yDSN8bE5jsXHVBTYYIZQnqBctLiBqgslYL90VezU3dE9kjR50Eux8GlVjad8gb+Bx
jIFi/WEYsAmUU9FlR3S0RlUd8zL4flSPU0RkgS15Cq/XmfSHQDfjKOtMhxwC1xokHWo6X9AHARPv
dXKipIodk1COfnVp+8iMRSHJj4TofohuXB+Nlf+L9nL4HHBE5OiaJ+57cJGa6/L362Kyhc0q7TWo
CwpeIBz2In1r0Jbhwl7grMBZ+GKsMXFjPWF8C+9o6Mnq9IBFRRiKYsPEynjktXBKQ2OUZbVakS1+
zqTBos6KOuymwqT2iTCXJK7Lw6qObVTDhJmSbwM9040KoVbUSw6xDaNjgpsSGPWWAzKIpObcT+yc
0KCUug5E8gFNwtQ4qhDdIbu8H6oQvAzrD8aZmT7tBA1oNqkF8R69MjvGs9Dzf93sQK6UXUN2alS0
GZigsc9r7nwsSIvWMVUU7bD+uKsC7j4NTojVLdvq3QnD2IBmNSO4/qV69imEwDJUMXDKJjqDrlNE
azZGQxX/OSnTp259EjrkFWFDdhcde/gJAya4VNs9mp/MfiVh+kq/L3EIi5FZbezHUeRk2dPqgfuA
HpkqCrjAKqdu5C6rmfrjEaGjuoXlR4Wcrw7/+77afI9jCwejodSiyhBmF8m+j1ImtE65F+1H/Up8
E6HEGuTkakHbvUoaNAbl7XkMrEBujDn8gfN7z8TlMcam0456r1S6BqMM8L+QF7CsLiXSX1e+EjvX
2S3h9Na+mhk2+BJLJ9yZ2Xie75KrikHL2yqO9sZG5S/jLwiukBGbZtDdvXgDmzzJ0BA8iqamM5x+
SjGJ2x3/RtDfGqT+rpUofruwjz4rkxxudcT5LkZ4cqT8WhOwSCYaLCpXhq510+bT5T9rZcqLJzdF
ptrE66plvxvOIp7ZXXWC6vcnQCjtv5DK0+vH5O0+sLoCWVS0OOX1XpA6thAZnddQppCbIFb1z0QZ
9ZVnNqDtDQH7LDnu4AN711kqESg1txpAx9F91YG+I44u5Stin+P6HEn/07SSOEeKeDiwqXQpqTOd
KL5hPYn+w4g1BEFcP8HNWQhxeVOqoJGAo5tpe3ASKLZEq9PjbHizSZnZLqYeGrFYnl+bXNqOU+6G
ig49JT642agxtGVbAGkpUNHrGy5tKt7ri17FKhbUBJ5W8fLdR/iCdL5d9ylly/eWw4nG11zD6Gbj
tvgxoWKgoLqNdiYS7FYHLJEFljZ9qmz1LMmbXcDOhllqnvP5ntlxtlstVc4J8mZrGLQ1FxEuLYPz
/hjzmXo2MME9+pmScw3FQPaP8dv8VhTQqRZjkdCiM/fi6rixySJ9etuM7mFSoLVdqWL1kr09y7sd
j7nx54sHZjTBdUy3xWBsO51Hw8stOAHt9p07N7Xn2XQWf9rhiptefgfVDYsSNAfP9JBxVpbKCOmT
Nt6ugNSMGBgPXZyn+VH8chR3auIATJudsenVBLfnbJvBXJ3HUVab09jM2NT6whJivHde4ZTQw/9e
0gy6+gGpqLaL9Sk0fSoB0QUxd7AzmrTdK3F+CYHJiTNrxM24BvIFkoER8yTrJt8HfflbjCHrBPFC
Lp7dBjI6e8922H8t6nAsUCD9Kl77kCswMC2IlnmTPZHUCg3zolIdvcLZMkiA6Hev+E3ONk0SMrcH
s1+oYgixdK1i2CpcATAAFOxJcHPZm8bEBYSlcm/fNAP5+bIjXpO1QzdsoRGocWqxb6TKtfZxyFRb
ZO+j6tbERZfkd3XvFezHLPBNMKaJt7cSWnCvC5L3aPwx65cEPRv5u0EfnFfL/VSHHShTNgFRpk4e
oOG3idD5xh/xnrptBE6LjTttzzl1p/znOmV8kxgua/L1MYidPFqQAX/FFT764JS0Dvj4Ad+o5ihW
KKhIxf+rKsp7QCIj2vGxJhkM4nRsLo/VSx93o3vjh23G1zaTCny0kYASDIr80zyFWaN8sVcITaJq
LYCn+GsWdrbNErwehyQ+UMFkgqjS+9WNq7+1rcBgCj6Qaus3S9uWomPaSeIhn9siEsgzLBFpB3mY
7iWjSX/wu/xX4sldF2aX2bnX8tnlGHp+yebQY0UTtVc5Bawm67lGIX9GLHW0qwV1gPVGwBK4rD8T
w0IxTFZYKDDvFdnUm4rioV7cxuj5wRJM2842YKvcshOjGtgAvBJiWcpph5gJyeRG2eUTfw8+nspn
gICQEkOmHm6VKKT0YRywBZgC4zRHGabvxeXviH/wy1i9HHZ03rGY3ltTSVGJk6BXLJWoNtMaJkZ+
NyV/aEQg9nzNuxTJKyX4+Hs+G4TsTDxm5Ta2j1wIvQdLuMbt77KfgPLHXILy6sR2oy+wPn456XuK
K+IHpck/1ugT295O5ceusfx/epkrTxP9Q+Ba/3oCXgydZ81/QF4aIb2dtsBfX1KPYntaUtSlyNFm
wce1zuWwmBcj0HaGV+x2ckPV94YNvkhjAmckhuQaci1QhgU1ruW0pSFGPEK2RqqT25FfcuPF0SgJ
jF+HFPSuvniko6EN2g7tdq/T2JsbMmIZqUmkHUH6Dk0SgEE0IXwq9mgCzco8blpm4riRSKzPpHMu
zckyFQVEG9GwoZnd09i8dwTfcou7llLiUL3CWV4Qb+2gt5HNH6Mqt37+uHggv8LOPuDIQM7DP6+h
04ft0+oynf4T4xmvfrT9i0ykm1K93s3TZneRkIa4dLlDGyjqSbobjwHMGx1p8M+J058idEJRyPq7
ZZNsOLoHzAsSx10luzyALYShnm5UIRw+tobuWPJQkDaCZee0fBQbWw5qyvCGIik9yFZV/p/1NafG
WxJsh9yC855UNkTdp897hTlNL2rHf+bQH9c1QimHYLcG42lVSX46cwXD3+V6s9UoNeEWA2DbtHAa
0udyqKM4lFfVnBXcnGrbpwxexDtD6IujE6XpXg/xM2YjwKm6DDBgufVpIyAdTPwDbSn6Qy0+YP59
JXJYe+bTHZEyxgjuQ7edYkiOeViGZYTc6tPBOYjk1Zy1s3BlXYrjl63EiyzS/4DAyg8nwyG6hxqP
BG56ZC8p7+tAFsLu5N22l7Y7HdfccolvnIkgFiaK9y9G0GOtcVcZrkvV7G7Ir4O/MYQ6KyqeaTOp
WW/MNnGf7aIUTykzK+rAWfznlXbwL787IGxw6rgYkolbjFXHl67GKclyIgHAk3tTLdLRz99LUz1H
0rxNCI8sZd8a4ZRqho9j36QFis7IpEKz0+NLzY06+wYuRsrgSGmcLQGHxs3jNhMOTc+HNZD40IkL
GF69HDe+NqoxkH1h5JRWMVP93e7HBsCIxU1xWwEcksASLSdEr5ad1YuiEWvtoX/IUBKGEP0PUNhu
ga+dIoiUhXV53Whxg4V6pLUpgqSjpmoVYFxyoFfLoNqXHWQiX4ZSsgGcKjHIPgiAP43/BJxDyCKU
YLIceWY0gFOruCQzZPfHUSj0iO6sxzTRLXH0fmZEiPWegYsvKHTEJRkDPGcckJJNwiDQ913WzoGV
bVW8UeOg8XVu506dVrvAXERdXfqYmFKfJ/i8pejWI0UW3hK1uOpi8U2vacoDr6IyzPcQTe9ct3an
JsDRGiniSD9HXQGy8MJ2Lhz+9s8hvKXwVe1Rve/hrhgBG1Hl79lh/15RmQKyvCfzLBfH1XvMwcLg
C1bb9/UukHfHIyGyhqnUumNTijg1Fj20k0SMlAI4RPxWxshVARyZlgV9sfYZtVVQS4UTPOZ70RQf
wceclJmjmJpcEgdxvqfy/h3iPsf+zFdDVj6EkS9Uqnf91DRHHJjccUrVnJRUlhHZihnayKaLukTd
dbD5G3tiuFTsS9D2TInIQ+H5d47yrc2CCyF1IOUQhLl/tvkkaFD7Tym9h4gOUQcX4Q1aEg9YdUMA
FXN7imG26i+UJAGYR5dZswnbqIA36r1Ucig2O7NoqNx8V7LLnOrUSbbW8jvUXbHt3JhtrzodIUIY
sdr+qM4VaWDoqg79o0X0nuIDHjxjv7JMi8lg7ARbmzTp53XzWkAJzdcCSF9qZNvp86GH9GTShMKH
EFeOXfZbsjLCxTGHzTgH+fkQzMTUhJxIfNxev5J4UkiGbKYTlDA9nXeKCC5rx003gGaWkPFGgNGH
S8+erJ/ZKZGeFvYjW+CZuMaJ7s6Zkgn+YQlXtzZ4Cn/iWy6zbn4Tbz9TAQF95c9W41ttrS37sVvx
1b9YQIL2cZXsZ0TmyXHkUvxFD4z+ekISXKKNoZ349VEXH+eTS2h28VwKyNIaf2K1i7aKfI4gJvRp
Y4YSOLNTDWnBrjb+jdQCkriIMeTSfty3biHsX6og1Wre6CYgjv2mWYnEQ1YmPNUISUVstlBMpVe8
7FbYMNw+LK3oaQu3mAlr0h7fOWq259aG3LLe5RHyQmDRZOw8s3/vcGfEzruOR4aaL1W+2o2GjOLB
dilPTYRNiDR0O3wnbaYLkc6t32I2PbboxJB32NsfjfQDuKlSRBvFapOea6/O5jmCGEC7U4rpGBdn
SqKJlO7C+kcryNc2X9UxiMbuDU5Fr8X1MinJD+RJlYXKlj9/np9NMAkDSYqRAxXRaDzSOW4rS8C3
n45A8TZwJw3xKFrQKN4tsT6QE+rzmfoRIsDlSksJvL4Vthv9zBPFNMtVeotTd4h35A571h9LmjXi
lMgJyzCPgFL/trX5lJnWw0Th1TxRKBI2tb1b0tHbJelrAlRrQ7NQ6nFgImCZtOBenTOUugD/x2Jr
kOIkPC320AmwzpnbJAZTeE1jIOOaNTJmqdo15W2qnvAUrNsPyXxEEggO1yo2M/TtQjHPEaz3q2QZ
PkWpcNKTzSsknsQ1T7YzWO86LPwx80ylibw/oLA14NoCvKWZvm8fI0BSgp6p1hQ7jix2uA/kEqe8
DU6WdliVb9HjVxZk647GrtMdynY9SyFz7UT6AiVSXAPyjiOIFC7O0rISseyh4jULdCasSaEWkSnU
14TAiAkGFm54fYSUXaiDuWgyvbLh6j83x9vjCY2cGU3esZSq8krZxbFgJ/Kw7RknSDfTTXrLqq4f
iehh6Ha2mNunxxi85lif77iRO6S1FPKsW3X9IaBbl0smhfUdc2sv4ZpGj3sAhdn7JBVRjx7DPSN0
dLvPrctdtQWTAvfA11QK3iQTJbaW27RjfY7sAWQhc9CkN0syq0g+u/dlGGkMSGy8EoVKI7Lw7btk
l7rAQhYYUIlB6mBUSwVNRc7kqtjd8bc1or6aMXMfjY2tcxQ/obFuWKZ/Qcswl33cvtTV6xl8W0oZ
M4vIHDDP7+JrgbHVPSHU8JRWsFCr+dLb54fgM/A3KNvNB3Zk3C+FVla/1VeGW9yDIfCwF0pDHUhf
FECdynVOsn5qUrXjQwTIT6hxcjz7Ll5LF5DjytSyAceOdyswyVedDotfw1Zaei42o6TGfSaaIhME
CYo/J7acSU28KSxsIQs/b6tc6vL8o/sFyHWAs3QQ/GvKcDzHdHOOgBL+jdLHsHEuZRoVe9frVybd
r5YmNhfhj3LAVSM2+n4N46cO/qDLfML4lyU7mG8FyP5Rc6rdkAKgXd6xntYXdm3g0KbIADR3Lv/L
0js4d+bPAd2l+L1tkb3MW6I8ZpSLY8Kobu0LfwLY7cplToX2kafVdQzeNU8VlqIOuO4urSBVExja
gPEZcTTyrsr/tmlt28O6LVMfMe6xnIezbQoo08uM+z1c0XhCwx1+g5DLyUUvpqwdFYOzI/K+GMrP
lRWLlqJf7HGfzZoYsWx7oHchypCcFpe/j52UCDtEtOo9oV/QD7bovgTD9JfXK81fuHxo23y9EiuI
rmT5Sjw08hngqsmuVYSDeYQeniPQVNCHUO1xNfaBBWdxmtdetuqZpG9L6/Z+oOknwsSHKRHki1no
J5xaTPW9C+GhAdSliZv3XaUSsg/Bq77rMPciymeGnBbZWdaqfh+leSkfymarrAhjJ5TAmz0rqrEC
hgmsS9w2FyiGgHREUDOCtoxgK8b6Za7wmWASCZq23BT2Hs3JdNBOKc6njcNdcQF8xwfCkJzTXtHs
2Te66rwD9Dt4i7pnWh94bOgiAXRadnCNzabu4/idEfHhS+az0zwl4XPfXZdYcmpdtis40SlYUSKh
xouvNzzb5KxPAbamju7mHM3wAf9yzKHf71BTEzggoc0zMz+p34e27hJkFPrFD+1OE+rTDb3oU/4f
SzSo+ykwrw7ThPpQwJMukpZgaYVRgcNtBysUZTY1cl5DQSxBUb4eIvYrt7TiOkJVZ8i7ks14PDN6
q+hhmknxkfyDJR8sMYdsBXPtG51r2uImW5sehpmnW/9H/UrhKaa1Fn0oUQcnxXSri/5A5egedXgb
MJTAWcw8X9yc+Tq6F8sywzcqELcwOuUwLFr/HqvlKwwYNe+1fU+gkJaQbG/MzN5ZMFpq08pn5WUt
MCtwsTVMyzBDcxQIFQhtFc9pVJCDVL16EeSx5HCWwE0aFW/MKcIiLHzTVICUJCAGvTzVV4lMUJZe
72oDIX6FcyNiaw3jDtqmAyFBDr0Ofccjb4rdjFQlfLRdXuvzTMx0oxn9ONMEiwmbz/SkBa4n1dLm
4cHtI9U3Hclm4J/gsRotHfXpgp94fhkURiIvII6Q5AJfHhPNyrH4B/NmRldkj8cwThFUrBD++6w8
tE+tl4FRxfQha4a+lxDQp//SdGKMT2akE8c9NdYJH5znlMayBSz18krb9poASfpJi5KperIDwuJw
4XjbDmxjQ16+dFB7AdjSgc93WaRDuuK3EGwRQK8y6XGvy+sWmAsyPfUn9y7sFJaJPwRsCpXwPNF+
B44OBQjrXAynhYxd6nwfkOLFIbWENdYbhMTxAZ4UkI8DIwgCLj745RH1AnJXoZImVxkfJ5Kx3mnh
3qW6aBwG5oOp5FE2gcwIW5KVYXIWkMskkuwVJHInT7nTlSJ6mCGEhTcy1pHqeCFT6j2LUX8zbJMS
pLtQjmZBWEalmixt+GKDgPKb4NQpFGvyxVk3ztg2r/FW2SV9vYxH1lh95BK98xr2Q8PT+yKTSCuM
vajApKBAX5mNoYoBZagHzl4EQYavutI1kYwovmAJNcY8fpAhUY3laGFs6MACVP6G7JvpSc/CGTm2
N98tgDb7rYpG/Er0/qBJ3BDpYnTCVa2EARPF/3JtZCddGh157jep7W5S/UnEje9YVO6E/jsRhhtb
S9mAvtpDcRh41+6GDuYQxRUFQp7cJSc/Fj1wlOlBqqnqJuTKfTaY0J7tT3719JaAW934FgArh6T/
S2z8WzX3tks83MZL5irN4+34SKmLz8DRkefvqFFooiVoiEXm1/G1HO2+cmvD4iIcxK+E5kcH+X51
7GNI31r3Hti2hxSe8Kj0BpXQ49/5pfftAdIhlfiHzfEos7IeDy1IVR4dc3ltFNPAJ9UCkL4yEd9p
TefiuF24TRB4gUdTC//zGYRIcRn3FaNrQvsI3WDDAGgZYaArfjZIUmWatBP5DaYgKCNwcgOSr/qL
N7lcDwVN5Zp/4igVtKZZspnP9tYzAVR0xTHvZvW+KNb6AxEYBgO/F/tYCpKyKMRY1iai1P5WJ3KR
+ccA2hSyqaWExENaF+dUUzxuRJEKV0iylI3heExKpEJMjefjB7q//C90ZMNELEfcIJG/88a64foa
sXJFWCeHN7i043a1GPSvfOFWaPhOWkh/b90+0Z/GB8z3AC5/Qg51OSAuOvuoZeEuNK0InVFiRDCA
W7Mx7kbm/BAzOacAfLZDYoMa/d8FPaJr3le4fef/bYEyR467/bf24Wq50eSpcW4uUhrcxZiWdirt
ZA1IZyCJidsGGEIEi730kJGSa6Qxg7R+55VRQmWFyDUunJV66am3NEbsJlpCX+v636Jhh8A0krIw
ZXEYQuM8qNcRAizI8/Nm8JxRhrmiZMChOMXBdNtdYw5xvkSh7+ffh31gxaPB5IrjDZZ8DveERgeR
epJmnoudGn3UiQgxRBz10bDqACnBT5Jis7Wj2/92jxpnOPqTyK9gHyk8ST8tPlVp3Ongwv4tBgXQ
tfsuG2idfXWM8OKivRCo6c3NENp64tSdomVdQS1sxxw/8M9HK+h9aIUu6tAMN75KmbfxpqaijDO/
CnI8kIBtSUGtU8w2z+geDcd5gwEf1hzta4I7tFibwvC7gjiQjw2wKUWkbkBJuILikjsEzi2jIlKl
xknxMOvk3NFbc525KM4Jc0qG9xuNYhx4Bp8AE6idPdRj76C9fNUbqtKHfCdrFpscc4IdXUTMK7ZO
55O+lYnF1HNyYlrjmNFQbybtuSqUwPWkDiclOltrjlbIR6PLfQdR5w+E3HcF5YJtB95PP9QLMmkA
kZGDvOUpleDUIsVD3fmohQ5xDQx3O2Wg4Awbo4zB7P1hI1NVM083PGpk+y4oxjCJkby5niUWKrK3
guB6zGWKiQ5//fRFm2ylDriZfoJo4lV3JYQ2FGEl0LuDUyOmwlgVHxpYdFUDQoXsskjMfUO9XNDl
LSOrtpMpnOnJrRokHQK37wnnWiq19PYh+se2+iKgdSrzY7WGQPwtvDbCEt3AoxqH1ZGuzpTJKNEx
5QwIfnXo4yNfPG/GA1o4DiJq8zBptcZY+g4nvr9L/a1iWNx75jKviYQ1zcIMX2Yqizu0XPn2rpDn
jEqLFwFWPUQEOoM6GD8rQvtkDTs89mKmfIIOSgrwKYomFrCiEJVCOQXbh4GscPCmnBdUMQg//w4X
8nxDS4DhU0qdxX+hVXcUu4PjoV+Fp6B92Dd9l83dbjIRXAZO86hFA54KTk+EtJtx+rzzWNsnpUJp
Tk3pI6ziyRmeTv3rBKuGKClXHHnv6ZuXoSLntNgDacEviYG7SxjhIqGZyLUzH2Q04u2ng6VZaMrb
Tkk7RFNEHAFTEouv0jT6Qd9tzdvsbIsLAiHvcg8M4MPVG8OkZhMWJLNcRah3mc/MHCuK6JFeUcmV
wNim/WTOxhR62KspbPx3vDoovRpX281kSyfh0LuuVIhHn1LUy6wsKeA8hxNP+Gc53NK42oVNcqe8
hBLpBkI74GuyZmrP5uOU1lkSnHbIXwfBIxgQaShwT431Z1MDsJJOPhdciQ4HjDuFyCpBLbM17TON
lp0T6nwT3Zx5PotSHFOnCxAYJkKGeKyIi8fiLFqaIlcqiu1Ed6nFrwPIRAEjRUytW64Bi8ptOdSW
pJhRJI46zP4a1KtANelPPui4WNFKgZgQcHtF8JWZl6NVmfk0JoZ5aAwp1BcNUmn13S56uKOeDo9f
DmOrJpFOveIj7ZHPHRjq/6RFxHjHnDkfNS3Mp9z5YDYAMvi9N5hS+FRn+8bvnjoPC8rzYWN9Ve5V
uLzuy8goeo68AfnT+DtU4DVNe90LkdwyFRanWSgDxxC4dRpjLsh/rhR3gYwPI2Bxnsw+1MjEEzzm
B1eqtYz8qonFXjkqyjjtDrVZC3HE1z+AVNr7DNH9jI540HutSUYofMu5H7gQ36lmno91+mU9gPFC
XipT0XdyBKWzQQDp+EUmX3V0nmsYIqsIZTQJ3mTHFQCIxQeJLM54BEoUHkMywkwZQsFKvEnnn+25
4IGeuMAnKqshE3nZyVtq7yIsE48b6UyUwWAYti7PFMHbIC1FXaGB/KFQpZ9bXCpcF+ddpTcPwhVf
a8R+qSKnbUX8MvW3mm4EuvmeNshtRA8hNUjU7Hlr8WcfHLu4D+BAYLH8OE+5541fhky1hMwSl84J
IkpGiLrTeycv51xezdRudcEZYCpRi2kSD+HLkaoBe+NZt7zDx5re9sAPmZ9S+3YkZ25RM+9humtl
s3MVYWkNwEJ0aaYHqSal8xrIxn0vIzqaDPpOROnuyoQ36fr6yyrAIa7USJKQK0034nHHwJPHspVz
7IS+5nj5wy0IDlz+3SmrSfNCjvrkFhR07xp7M/uDn/T3oJLmoJxOlpiVmVH1l/PGUVfPlLERvnDp
20iAuGj5J8oiJGibWwsAPguClXTqP9dIytNvHqDQUV1b5VLQuLri9rzv0g7drTS3SGyqOAqg+55i
R0ujR8kjIhrfdatjgBDz1R7wz4SmhlQd9VDzFyLcIAt7ns4pnTAcpfDL5n29pXP5te56Eavx60AB
3Vd1W1NUdWt4mlRqN3Cff4BBmwMgmiuAVHZDL6FsiVNytlrtVojC+i1y8KbLZXB00iO4plbTzOGq
Ic58bYo2qckTyK0RBgLkvD/zPQ8aPPmimrs2GUrocf8z4H+WCWz0aULYcI/Yw4KSnDA5bumOncqU
tvy6fjy7l417yIvRU2uqtfvSRGvk4QZ4OGcZLk2KK+44/If92ZD6a59wI7TU4OVsab5KixT+sPgl
YWpInnqbo7NdD/tqdhR75XAkM0Gg+abku8SnwJ54IlECrFCTXsyB11EIVVrFTun8UP6IV0TBrJuT
wr53bme8Dj0cwO9d6UwDKwW7J46OyOgPp5yvtJv5K2h23mFNmhS0ajRw7JYNnbIzrvOTWS32wrGI
j1NoUzr/4Dy+drC5G235A/YabIHn+VMqYCCjRTkWzFNerJyYMqgzdyH4jomxNXAzhlulC0PpS8jm
m27ma4L/0WvcuTQCHQSt+FITab5lh4yZPQllbDVxJC/tvT8Wf99WGu6Ag0hEF2qeZZi5p4XQkLTm
hjGbnicpSZUeLtnlxmPlfd2alqMsz4OGTjCp3Q/4ynliGDeKNeOoHSMKCpxXfeEhpJVDXHs3xqBT
ddxgIKafuKkKq/Svw0HHGeTcpz8Hsq37HjLOoyklDDocyg60j35sdzlQ/FGTbaJwMAbAEpzv6a+L
evnavRMOWwAs4DTqdQZeY4d5H0V4nN0qYSIdUFCd5Ftmk431QzSZTjJzHrCdJITJy+WB1E6YXW8Z
L+m8WEW6Mp6f5XKCofsGose0NEqEQhWljGCA3uNeWMFLgOIts881SLVXQM+aEGM2z0YQeYalf09f
39tyI5Yv1ow+C4FbGGAYCj5wiRe45jPECu26iHWy7d9VMbg8f3g8HGwfe+cj1xq0X7iQSrJrWx6i
sHyww9ga7Qq/gY4f+3tC7P+c51+j32H9zIovi996fozLgT9pvx9huI0J2Sfv/dF1+QtunHuqZRpz
yK/zaWaC6G8rPUlUBymHw17U7EAEom0/USmZ8BXsMCWxPgasrzv73O+SY9u/1dRx1XOZe3r1BFqU
qeq3lzFEy1nh+pcQ72JEx5CnbMrYQRF300imi9YixSsyceuQ1jx8JjJTyN2zLOdXXPk0iGGfF2MU
uP1Xk8UFvfglyTU3XBeTSjxrcI/EwUpsCPgcPoUVmbnJDuWXhQxUgoZjHdDWy6xjDJ4TcQJ67Q59
CZE8sDiEPwyF/S0D0O3FgA/9LkG/Yue8svyoE5aegji9xRGrA5gKaGM5TZJdsvayrUtzCeN6czMz
ELqNgiCFAny6/WSnRAreFhGu3C8/YxR+sxvDopwJHGXZUkiNtACPMBfJZVTDs6vDlfdbrEjiQrwb
k0a8tb6qfyH5jC5wbZ3DsolsJ5SGzp78k3ADILCjlSd82omk/KGRn9qWbQ8PgA7V1pUcAeR4TEnR
G5OBaECsvys8axpB9gWZ75TTPwftjkA5FPgo46IOGZwW1qn7wS4DYJh+v0d59MS9NxbIM4n/NgLt
hWPZf/5r51CBgpKpV/2FMr92Ocs6q1exiTg4EZxJ3q97CRtOdu5htaplOnHC1qTKUMnTrGJXaBuX
1kDHPwLwSCjAUvHM6TJEZDLejYu7Fg22lYPBQe9NRJA45PePPrjeFI7nF1IiiQeTkzyzmixUwlU3
D+Yk7cQ9AJanZ+6IYTU9naoFJUwV6jKiZTSrPEud2oQkX+Lihqt3JGA5pYbaPyzTMX5z0bzM1IH1
5AGHY5Pr5UvpZqytcuA9oNEdqzwmg5V8QznThkFSbP+rcwHt3woVthp/hIEIfr7zT8AhCviKokqX
uscIuQ3NKrstZ78jSOfs8BcvqsJxhfrHvqE8NByOoLGqwGcXfvany77fcnZzLMGd1W4v8hP8qfaa
2rFWtTGblo/291OTIrpYBnIs3sTVrWBbNPgfjLd13AyHEnIC2IwsN25WXOKjufKtXnTCyJeilYFe
+nUOOQ+f7ll+wabtaKCqtr2k7+Hwep3nBLuF9NuUSu99zs/GG5KwegHWVZXgLAdDQy1rIdSA9GY2
+q/Uu/h8hQ91CSka0NNeN1gOSPSPXvJuJTwRILUe0zU866paNtINoxSp8VWhdV2le3v4XIKYqr3A
JOLqhcKenadwPtg/qWD/63o4Dev8CIkKmX4p3oGqW/qN3/RXSgwmjMxyKye+DjDDk2brnzeJaHgM
K7PLFTDDJw4w1PyqfykV8xHqg8mjBb5+yizNvoSQTSoCqQGDLFz0SJNli1/YeHyC5q8sjoBlgev2
4LhSWyYVKBRw7XJ29GdlwmxkOgVgwcrKfBtWMYZBgHsxxNbTlxobpBRESfPhdgAzoRvG7TtPrM65
nDDRePXofif5vlOHx4NAJzB7IdNuhvNvP4usN3WFKHHY3994KGIun0oiIbhTZedVWAY6qeIdX/Mf
K2gk9LAAf5QaPD6oNPyi8bh0ZyHKrZhLAOC07I3wyoxeXbLtc3CrR7ezXlyWwmAvAtcHyPLETEzV
pVgnbilZhwHEk3oIRcdsmoYP/lvYeVNahqydbx750Hg3f0XZSctr7EM0CrTpYYU4av++7K7jJSTw
X8YpMIFTyxPQZhqNXLN5K33LzsjJVBG0NKix25caAtuQ/4jZ5gcWUOBVMqX2c38cWmD5ixqARfzS
Plmz+wvMYp1NZUmvDPgti/6ss2AVnvVzFsF3PybuNygh5bCMNsfpcmR5Dqx3PdVjgWMGFlxbR1LD
DZIhJg740rEdPZUOCj0LTh5AjsP/urlbxxrhFgJUPN6kLr5IAm8Cx1DCVVrkoKz5w+TLEVpxCAxt
VpKAbfCGKqfET+O6ZGP2KbLWXhy1bZAkSjqrrbZpb7HOEvJi4PF5XCbmiEja6LGgTl92TmY9OXEf
rNqD/jkoreISW8Xm79WhbPciVPQFgIfA36ZAupOScgrH7oDs/tVnQMW5TchG0xJSurWsp1YRx7/N
ovGvOZfP9lN7ss7xf4Gunf+PG9hFfSNv4IXwZuH6UpNDJlBzSrMkRA3p8aWTgnhOutJFa6RQPtiL
o0AQENKOQ7cDB84KcIYMBjb8kwsUtZB/1iPEMsZQ0uDETI30DOqM59UoGku69r1N/E3KfuQJOhxl
9QPxKabvp5+6hG8Nvf6CKOYVDBkzOURtCJpgEOIjMfX/MSBoCn1IeRR07+ZZxDYDEkFJ2OnGoKL7
88MbkBR5jsW/JK/6GqeTGpvfphUOV77UMOuNKKctdFVYIv3p269xlljk4491yMDRwScR9y7/CXDY
4F85OpLytWudNF+DJ9WPGZi/MC6TQ1diMjps+tlQi/t53RYq1LktgWhZ/DoMrS9Rd3DzK49JIlhP
8J56HXKBcMa5M4orP61UCx8z1loJHk6guBZ1WTzMe8xMjRAPOY/ibjVwLKF3Q49MtaMaTqgQ87Vp
CcN6A/upMCXhcfycgmTMOsz6cqgsoeoGbFXojeCgk8PEASAqEcdaQZsWn0u1FIGgMhP0twCGiDBc
Vh6POZDoCzy2+RM51zhFSBc/H47h0t92AfuI1o2cLD3NGXyZZgwW+SxX11zDimdpT21IRcC2i1xh
D01Fm1MxWuujiQ9aK8fQlfeyfwNZySXBVST3YMzCqsLJGcQ7JHl2AGd3jJKW5DIpww2536cI9Zbz
ZhdGsX0YIlPZV9MyOG8Rd0iEjiuOZMaQlK5NN2xS7sLJ3Hrczhj54rEGFeJjjlmndaHGfwcZCBfi
6qiTLBZ0HshIz/ZgiavNS6A6af+F+XNZjxqnCxeHbwfl618nHEg2cz/Ddn331nKdFRsaeCvdjpAl
XQjHifEeO0IH1/Wt2+DLD6x49l6qVn24aakcyVS6m6CPgDCKAp8IwImiNs5PdOTdBjsjVGpqIBoV
A2DEBxpMSP0bS6nJkzOGFncEm+Hh9xCc5nnY2X4AJ1UyJjxL9sEFtTUzYUcMSEvUb2h4H9DAceQZ
2TZ4rv//K+/GeCBinSleRTYT8rwbGKvz+xXvBHsKQsTtnhslqZ4Vj0Tum7i4Qg3o7C+O+HUHl01M
G2Aac23sBP/evHAXeYLDCVKE5dKuC9tQyOxkZpAV6sqsLXYRkoiW6FWNf4GI/0j7fO7Yo1WsdxvS
CGjFDry4vip2DUMmpem/1KnFFl3/VteLeUv53TL5cCHnx4gbu2fhe79Wgi5zaXF+0wc8dIA4JDS5
vVV0ztoe+nOgUB6+duBdF4yGtm+Kj98XF9un/AiaRbZJs/ZQAbTDe+x1z5+cp+gbqa2FDWatKVaG
QmKtsqPmK4a5yEOS68BcNUEiezDKxuWnpyAo7gM6+wRdJUcmqo9WoPNK+hAH0za1V6vYpHZr1KRv
P8jfCWNwVzHx6dV5Ib6MGzpTCnqkcX8LRBj0tLpjwGGf2gqL5nd9XtLj/u6QGQz0ldP/YwUd10KU
VVtEkYO3mVomUg88bKHvhlh0AX97T0orf3BuVyAyico37EfLFVdRjJVbe+RdU3zAapfRTS8QlLX9
ZvO1cZ7m7sF9eJhTbg/B9ohf07O2tLF1R/H7Y5taC/WG/4b73pIL5K4Esh2ovA2H8sieyWAXCTwi
yBZcDuLCY8gF//0PqaijRVtZDm1zHzr08+JnJTHt1bYtCaRx2nw5O7ORlODzo9FMuMQg4Ca27pBv
yNJdXFkLi53ZZwY03rC5n3CVcJHZuQj7MtGDsLnrC9OA2JE+wK5puxj+t7I01hFPJO0igQW1LSNz
wj4SVH6UTzfok/+dSm5vZLTBAtEaWkadgyie269Tsxk89wXidLGJNzgNaMNck4WQbkVEvV+Ty8Zy
HxTuQCVddQSeru3BQh0dS/0XgtQIUUGNDDtL3HEiWHb6pJsQXax0hXheVFbVZNfN1EQagG3vZs9J
aR6IVSkVTfkq3D49clLev34ZWlLLOiZLX4TA9y+aZMjRSyfXeRDEPpLUy/iBaG/uhSxdvNNd96fU
DsLDI3A7mfA2C3KzUCouV3ycEU2TtazTa52hj0y3nDo8YBz3GLrgDvl1bVaTsSVMYmLZ54qlTkg+
sqGk1HsxV4bR612IBhBm0c3Se4ly9tnWC7c42YhwQBLxjHi0C0cHA+V4uXC8mYT3uVcRLe3B7dXU
KBNqZwdIrueihYrkbuXdoIHd14RjfBJsrtJgQzLECEUGIEYvocbEM3CCBoGSd8wylDkjQCXz7K7W
MPF9Hf4nRe8ERin+qKISksXHPH4l6F3Kjf7hXBxPkKAADoizW0x7mAlQ4rTxh44t/1tuBdu49iVs
3k/Xdj7sWJ7Cui9aLfsdpcE4GMEX3ksmrIxYYjZ3wmRql373RZcSgNcNn1SNgDFbu6jtLHyZBlTi
TfkdAYZWd/FRxF5jdxvPabcV3sNUYdYm3ZKQFnLTrDif7UGJEH5TD3+li2j5DaWDrhbbFC8AMqEf
+tfbvsEdVB6YEBeJjTBLgJ9HB8Tlu+Z8V75/hPZGNceGTaBk5HOEQa/34fywy9g7BVXQmoYd43RP
C12LZrLGDCCopvanD5Hap//YDxPUqBAKmjyXTHl8feStvrxEC9l/pG3RsYhyLJjj2Y/prv4RjU7r
50omkGiraQq+R+nyvq/OoyVAuM2ROTlQI/Fp0EftOPu0lYpvAQgJ6IPgmZdVjOgrx0DIcwJl6fx2
wCfFhFAg8PcBVYhZKImamV8s9lLCFuLeXDbWmhTYH0h27/dADNfH5w5Zvmm7ZLLvqCquHWO86Wu9
ZlDkwN6qcjwLKyZOkY0GysTBGGoyTSe5xH2rItSGE0CptiQxfMx33TVoC/NX4sqKEvI2tAj65jqq
M7CeiUO+rt6vJEyHGpHqlTw6PyySOoy4jzdSwFecTuz+Sn90ni1DbUH1WJuFH1TDn3wY4DKVLltz
Dxw0ND3DlBYnCrK1GTl6JKi2aQ4NDsspAdp51O794cOwM3BC0tvmV7/kp/klRVYvLUVrTr+jWyNA
gUab/RaSSfasKsk3rXJZPw/zCEExgvtBsXjkiGMTD2q0OLCPCw17qJEmEOeheweKZBmlmHP1UKhL
iVUKIe+gubrwuZysC/b2DW7/dvuFyYSklFpaCv22ScIPrImWhNzjQjvEBM/iPfj0Zv6I64zBb/9v
a8SzSCqz/ZguGzq97NwRgEiCDu3+IH4XwVhuIesGVp3FKhGlXPSXFrZoYatYkQ8xxJSTEnrcBiY1
LNspAurHRpVeOOh7LwPI8P6aUEOQCLzPAVCkkrUZtDCiyIhkbnzKnsTdkFwyWOeKaW/4KR9A/CPZ
Wl89EJSFfA+VwVuo/uOFTltgo5rkWvg7+wq+W0D9KBlS2NQ+BjJcrLOv//gZDH1VHFssGeZ/LA8/
Q6TTI1GbPS3QoYoj/AitFTxnUgk73whkH71MnYdQQT9n7+GKPVcc4iAPcof6d7TUR78fmPu2uOtu
V9uxSiOnf/Kw6l5QLDfezgwZ8sz9o7AjRYcDkL8y+fw+1p3OzQH06g55IMQj6/Yr+VYShJlyfehh
1nAW1i7BqDyJ7DSkHB8viMmcsGpwHyFIY4RdaSv3+8DYcCKKnm2BFI7OeYLwiKHY7P4tQFxPOzAw
eoemCbUiMLYuG7MW+RVR1rQqqV65NCTwOrzoRFZSCUungsfrx07Gk9jZyaVa0brRu4yvHoISbN1B
XIb4ID/X2HdUxaSt4sXWpyhpcafeO64ZJX2K9FnRO90xOoEDzlvwaQ+Bfg+PIq/ZAM06NoQg1G/p
KHa9OeQl330cf/MJlClnfIlKI697w/p413Z8W16fBMDZ84MhYOf3p3Fn2vGErnc7RTrY4Ykr/IX/
YRwx+tk5YR36r0tr5QxIW5pk0RIATuQSVo8o+0OlmxBPtoO2wnjSQkIxmdx35FKH7t2fFiOxmdYv
l99eebUTPo/602GzO6l3nVQAvSZ0acMaYrkr7jt8AZmxy+dDX6l8drMwh0c5/YUlQo+/rMUCxF8R
9tGdR6yGM/ZIJ6hQC5FLF/qolimhDA8lb4mK7yUbEIF9OXruZnp2/LfG8RzSYnzTq/0vO3/KH/0D
9dLOwCkgBanraLx/FzkcJuf3WAXe1PRBf8qPj1MJKT6PHMndYna+eivfWZ3IrmIHM8gk7SS0JLP6
+Al08Dv2smbYmDkFqZ44+bbGl8cDKKuVHe4fHSF7P9jhpY+QV/Y4X2k+G9B7mUZa6lZzPC3aU2ym
63NOjH9j4k6rNa73CPYm82wWYuBut3JUo0uAiyqYNwjN2AWTleopefxVPw2Elj10RVkFmsrjoyZy
w8XDgRGbob417GHvLXNr+2EKY9+/9kZ03qgtceABIpUB6n4pe+mMhSNGyyrMAMvxQr/oQhXpAZlq
9AGMCBl3MtuC4Ptojv00CZX/QolJbz4T2UKzb5T1wiiCA12PYkGPd7QfAaR3Gt40I/P386WLtWvJ
gLgWk1WLbj4UXVD5ITaYBFvtIbwmlmdglEd7u2MQRDa/PxSYRT0uYEQgFgkd4CQ/SYHO6DjkdHxE
vJ16SgSxtOH8KSN+HsgtSu8kfAPGGqLOjJi8bH56EcbO/TSLvrFJEPCpN9GyngUoKnFrAgpWNmbh
u3EZP8/t+ifQJY/eH4QsslHsM9+I6+DVuLb78zS499FKG+RxvUOlVZqCOmToaRfT4KU1wmn8+WLk
KIXg8J+lGlutPZQKfaeTCmYlaB+UaKW9GzWhttQnD7vzuNKQMeS/M9vsN7bjEDPmPbNze2Z+pVqp
xAsOsHiUIs7EAQgH3EmmKkUJ1KhnR0ewAHphIpx7ryKAwStHnk2mMsBUBEdN2TExRSjF4w2bdqAt
jof/+D4EVbjipQAf8AulAZz0Xq1uxqEsu8eQ0pUARDMp2L6wfUas+/mlQmmWx9lr6YUVyZ7b77//
5fl8M2EmhJ3SC86ghlMU1qstJzIfzYoOEt3uzqN9cqdELbomvo6HPJuQ83k5DOQRXNYCFdPe4PiW
xhUyQ3lqh5ufg/MRmIjagoxgBqNiEND92LPv2xDZ5x/ygFvSurYiZj/ht474BDqj0EkaFYM3x8OQ
2FkAiEkXMGHrol4G3ZPhVn63AMN1oVuHweGDIZME0mTZrd1h2pr7IGoUIp0YjVAfw8brwXZNgt8m
skzkCJ0kzYLnFlzwoACLivdEuOEeLMOtCg8dEY5g6k+xKu6j3fschvvyNHpxYOd/9yZylxK7LDiC
7DnrsCYiAqjxn/EJtQrtY3lV5QBEL+1gIrTFqq0MNC73moohOB/T2Zsv6cNbWQdRPD4XsWQ3CFZm
Z3XM7Cy+ync/8H3M95jitG90Eu2Ml04G+JZUTM1WypnjTQSLjBinuXerSvHlhRdNndLXKyCs099I
UjqZFP0xIlzBKmu1dzFcNMQl9bzMZnQIc7m+NFqyo4AtyiaQivQ+IU3do4/PpkhD9DaEdXefbgEm
02I/gwdWVQ9GnRcCXRguh2sud8hzR+hwIXtamhi+KOs865ZQEn0loBQ3t3fyU8oo35lWxBOhFQdU
nTKM93WwlsvfbzNwdyJ+Hx+NmITUwg1VvAyhPM1uOErchyQjjGEYYC6a3Xlk31k7PUs7uHHlDuLb
9lOwmJwUsj5rq/rYoAKRKauSj4N8QR5xxOT6I/UhWqPDrClMFtweCxPmDfbgwpkHx2yF6CqTtG+B
zdHkAhMlYhLAPKJCybAPuxfn1KVEiRnzn7oXiuevHqpohM59M2Jj6oF+U1Y+ba4iSGyxaKOl8/BY
jHQrgvsHQCyOXUtiLtX1WsjnbLU1l/ugQhWm/8PP/vf1qZdVBpYz21tM85pPSNrPPkEim0U4PJIO
vraSPusxrfK45njB5hlrc9INWEXy3RqDUI/f1TA8X3EVQkOEK/VlNzv+G7yoq39DOlHj+ZgbX7iL
vYFC+b3QLvPNM5E/CofSz3TzJ2Vf+JRz2x8fPutGKLEJ3fwBh3HpgSeziFlikdxQl8yYNbPEz7yL
19I6eWF1jsZeOhRtKUyMHymfiMayAmoUW3bXPpQr5r2aTPIEwPA707EpFgHR+/jr11GvtzJPupa2
NtVcp1bVtpT9W8w0d1USLHWTRLCZL60XrtA/1lFMyaot3NpxKJhqVmYWgUpaOMWHEvGdgysOuAu9
iCLHD9kGmDQlFXXlzc2dEdcuJxJnwWfIJNYDzNCf03FP+SVnv0MaAEraXfVTAz6MLO4muRgyIfk5
qBz6K1EXG26N+Ic0umiQUV35PXbzvu6yJs1DRisBXGcq3/UFkF3pqKmZBYya3t6SgOIqzSC1SfF3
9L6Hu0R+0rRMn5sbPxFcTwNFKW4UWwUsZgy0qtawoGd6As7cutJ9rlL4LWL2EaFHs3+xy/yjN82U
Rchs3GlV3Xkr455xr+zO5yS+okrSz6z2vTCYWUH9wGb5q6w0VCOnQT9an3nUpXVq6gGCJQUBD9T8
ndgL/b80DN6eyBcLocPjlEg4hgtq38I4SwytIhtT2bqhQug0msTiLKSX2E8AiQ0Ws6U78EGEsFVa
E0iloCtGHDQK9iUgi8C7tac1zSm16KW9I7jltYTJQRrR8yKY9lVfPdLPXwxq1ad9q9eFY0uIGIxS
gfPnM5KnPkrgT7qE0ykoQG3g1xbaf2Ju1dweBTPN94QpJ2GEr70dP5k49uRMLpJJDt7OFpsStgPB
a0wpjAO4fUjKh/wzm4LtyTQZV7g/oP2bTAsY1sXCfAzutpvql0k6d3W7jPSQCGL3F3s/rDXbXQlZ
nwou9khrdwyKuUahoMbrfiz2bSMo5jITQzR8Ek7fZCimzUVycQHLa0CNeTm6FXTUppQRVwRUF7qw
x+KC2ZmiY6kuDM5cnMhL+m3ZhHjU6k949y0PwN7A1gd4tMvVk1gVxr7jXPuxLasaCwAogJObEDKV
1H2MYOH2JbUnCQJAflH3y1OlZCZlbTauH2jTYn1HeVvla0geyTdqg2klIECnP/aNkf9J91uFBgUl
X/DcX9SiODVwaUPIMTGpehxDsK+4KtMhrbex2kMSCpqdAPkUwKKtPwYI5oxk2Ortk2UF0BLyQ/E7
Op2OyWtZaw3STtHoP22hN7hVCqhUeOTOk/TXLPhrt+Z3a0FzMvMvBqDjqD8+BXRrpO0A2xUBLSdN
cZtZu5rQfah8bBN95HqzmTw8acrgh0fwlMoO/2TALO7eFdL4NSy9TIk8IZ8kQDjMw9jNsB3uvRkC
VfXZxVt2akmmaAAv3p8ifeERK6WlsQWMbaGRyWv7HQc2HuB+IhRoM+E6nkONlKbtlTGLqgyjokVJ
CuOsZCxzxQPePpKW22S2HBFk7uusLVlEJewb1AX5ra5Ffu8/gi1iq9I/qV3WrZzadvvPnj7RBXI4
zqE4hm4/tVQeHzyGnO0zEen82XfVKCPKCg6MLvC3WCTPnbbiDUFZVym98UO2BLcVjbbmwuc70GM8
sQC5XPs4X/ndvz7wIqFhrzIzS7juA0PqHT7z2ZTjO2HZtaD7EpHfly2B+sIgJn8Q2CP49PI4V6eM
1oLr2uojwjstw8Dzzq3O7b8+KPUAFeo0U0I/LK+z5z0eGExuE4Uh/elN+jzzASrP2s1/DQPDSu7a
nDY8jxxsSdlsi3bEtNzHn3V7v8yl9J0PZtdP9cKMFoQIg2NPi27bUcmVdy2we//MzfWGJ/t9DjsL
5xzJLQlEUyDY5OmKrhO2uWXnDTdPOYNu3ZGRh2S8hEG73dtKdMaL9c5NPSRL+N047XHCF5HKXuDN
Pk/4WGVl6l05HmJJzO0b2d6/LT81TuKJ9vZJ9HfQDQABpt6fhijFaWgJUQUS5rJ1p03VrvbLKLe0
BhiQ/FEx0DP02Jp/SFP7oOQOa92AYy+a6nDsNXKbuMcGK3Fa7yTHD+b/OQVWrbc/LYX4IlacnFkE
7PyFsy/dt/Pxo8Ex4w6cAGNpDG0FZh3DpcmZ2k+bHbJ9Ufkwigh6NuNrV3htmf0v7TRTadjhoCXb
fKGh2MTdBmXXuYEgiIxFzmse1v4iTg4vOnVROUvymRBiM2HruofaZrPahDjnDWTGp1lqEeTA+IoD
o6qhpKf4dgYUszMBVYsZl3f4IJ6h6QAtoG181u7BM7hbd9UgjQ2hfGmWeRBedozj7FXUlOpJGdum
l8Pi3ruQ2+0C3FpqUhcaGxIr1e7QoKTTnlDK8wzgbDQ6hkwBIVgL2MP64NBDxgyAWAkIrVSQETY6
w0DSCvzYFUKe3DyDx1+v/88mX3G7hLWs9sAAdD5I8jwzvgXv65FYq9Ai3OJ6ILkzrInrI2r65YtZ
380mNXRhBVVg/ZMgBNr+zTGeSE5m7KiE31F99uily7Z2/+4skx5d66s9+fHe+NhxW3ORj3hLgOZT
+ebZtELbT9b37pXmIWAhSQN6WAwLs7EZrbRhDOtpySUdXtWxmIMKosEc0ER+UfF6VemughgoX0r/
c70UWpUwz7gsvsYOszvu1Bj+mYhriWzO68yRIVcX52WXDBYlQ8g/RFVFZX6ljUrQh49SEu3wiru4
Vh4O12sf24NVerVpckfSrHUoOZgND0FF/OMttdOPWsW1498vlwLzwQvi9w8+rwc0mwBZvuCbG083
edcvie52blzsbrFvgjvrFXWUiIzmO4BoU4x1+tl6ZK97UMeiaW5Kth+v7OEBio1KUOayBBBcBL7s
eTgAlNrEau6ClENpxIqOMzU91ZP7AmyKHitZSmPdLjXlHnG+BbhaR1fyndmFZXGI9yB1kYx/+2tp
KWhs6dT65HhbKKLL1E9QyWdEQgjYn56z0j1ffrI4/91IMdrmjTGTFJ+8D7KPCtdv0zK+6HdYD0hv
y9MLpC9qayri6H60veoz+4mvwBc/CcenCJdk1YlOB1RIeTWhbiAot2z0t/lPIFUBD8cuAhUV9p5P
qIiQvYYdrCpBzKWgzKYN6Zje5FodslaMN2Z8TqdB1OILiSlTgAc/nTIbPeafpiNLWDSdpJizE17A
Sql5DBVHCzqSV8CIyRqW03TVCGXfZ9kSEPcdGIYML/4jUXbrytwMkR1tyVvO+7ptV2B46b24466H
MuqFtFWCcK/rmKBwF7qhLpo9lAm5M+COhfblUrjac7gmPQnFXJNDf7tfucZCtZndXg8ANkh2w4Iy
avomuHr7n+SI9Bu+DfDiN2xOS1E76l6JQaPXji6tKzCcX9C4Lw94CQv4DlowTsdLFPAgr3vyfDoN
roJJoA2JWd7sQcEP/O+fpg6gbvEJraxzLO8tVWiUcIBiCcTMURPr4+/wUD4VIS4Xs3ftmFMgQc+O
tMY4BtSXxUSLF5kdF+LrU1uLjxcmfF/Xxx3X+nVsnGJ9piudlpdanrXsXMfqF8gHPwm+gAeSzgxW
Y7pNmspUAuhIWNtslcYazrn9JweqdKQw0TywkFc49fKIz4sUaZGFr8RXi3tOGP63bjHBs7W4yaTf
BcVGwJZcMB4FWAnjwg328XnHN5l0ZYw3PYrzOPo4Kr6b5GSKrBDWYeQbfLxVzp9njt9DPLi0LGsM
rLx7gCrOKkuEx+JRcMaQE0hS4irmTQfOQovGzQQaiesnCdnuqzB9U4vNIiJUtAD41gu/jv9x0XLe
FVGfE/CPg8/6V2jPHH6q7MRluJjj2qM0iEUEbE0u+nX/ZaoY4SM1v57voIvPqG9PoQksQRQdTaGW
PjuZy6kL16xDnFUSPq6jbz2UQDq5qcj/mq8MiXNaYUJ8K5As4Cc4e3enkp11nZv1iVdc3IE11IYz
hxImdy6MSejvA0TNelcnTf3nnlzBJhEucLd2LJCQVL2/SB5JTzEZrAGv85ujMCNlmnL0IcJa9zBH
62lw5JwivQs+cIxtnn13h+tFcSb9zTEc+W+t6QzQ0UCrkQ8fzpmaAnQzGErAkHeF8Z0wVByYDP2e
5tdEicC7W4aAMw5MiTTdQxeMkxudY0MQf7O5aNMLoEowaKv/aebvtv/p3Xg5gKeS38C987YDnh3u
TwmGmZEXTvzjLpdQeHfzvYo0dTwOd7Ffzo6uuxSnmK35lF4cLLV+AT2rAacmjQ9XvjsHQ+RCr7di
4BwzZ8dtnUFep1laN5Y+2nY/IEzA6h7K1/E10zIxNWxCrOUpQC4vOS6Jt3cZ8PeIcjGAd5c8kMjf
euull9Mugp3bRCIIqcf7q1Yz/66YyiwPVu4GQmZCRbnJowhROz6QCidhhJwiSs9cykmXVIV9wdl3
2KPlM2I6iWKdRf9WGw521v9H8KBzFNsPodVhIejcZ/q2+1VBo3VrcDZNpGDwYoysfYS6rQPV0jqC
TdAtWv/VOvoe1ADMbkfqi9vPKTo7gyK6OQnF5ZHKZUagNqlXQgWVgvbGr8ztIJUpcy6pviCzRLUj
sspGnFpBsEOjVyMlholtkLtFztq36Ld2JNck/n/nperTL1OpncEDPz9tJtjO36d7BVemjfy7+0jn
y8m8JH6rEDzZ0S/YM4GPnbw/ucRqVuwtbmiuzkBKWIWzrDTq0zkKzjfXooiSl6Hz9HTx36Fo2/DI
2mRdzz6SXFOVM8vCtBYO2dLUjr6wsLviOlAVLoPcrZmpkrwz+358FUbeLto4XH2Shh2FV2CwGR6m
C9lod2niiPsMwEg3wiRV28zvriLSAGUW/Xwx/N/NABWLdE1HqEAp6i5U4lC1AqUbxWP0bFL69QDs
DvA+EHPanIsfBzipTAILhRpQN7QHwNkgE0+pQWvcWEtMi9HRS5uOJCkw9IcLMP0wSfZQmtSJzYGF
plblISJOKSmMCMqFTq+9itYVTr0def4nI+yBTyjktsjsVN8M3XfEl5ydmQRDrdcJ2vFcwWICopPJ
+VlDearH++Pq0aCEhvujbFUdS9mE+J/DX+SYi3nUw5F40X8J1v4GwqO6/EaYRUGYK5P5xtknPKIy
7aD6qbrDbvO/bkv0kOAVFu9nTAqtVTEXaEMUFZnIe1JuNzfVdTaetYROJsMyswgzTL/WF3sIVCoy
ebhprIcD915IZsbkeNxNI8RehVHmWbDq7G5i0X6lG35f2fhFc9J80RvRDr/AhBuzWdfrbNeykOFD
0WeNvHQEtCjH8Mq5NU9cp1j0uGOxlulCLooJqbcpqUFBw0OJ9x2XTFJ8ugW8hLGt5fkfG87caVIQ
dExjHoysjp9B8kuwzG9uf2WDVI5ObF93nqPARzfNSz/bODCjsdleFfinugZJGZD1SUi/NCbiA7hA
DRmuc+M/Ai47gIjOyg5bsA54zz6rqJoR+x1P7dI/D91SIqkaV7wErqXyIpR7O0cMCOVZKmMLkCV6
k4mnnPCNZk9Os1DPXGhQgLj++juYXZUNHwl9i0FQLVnUa/VyaSsWrKxx4Z+tlnwm1Em9NTiUGA5v
fcz2f3/wIMtO816+lix53njyoRddvjAHSi8CX6+2ZbSfxkWiMmkF2wLTTxE5Ti3r2RoCbAVgCCqC
NHZ49AvrAaGWMmK2yVOuIoU2StJ1Dn5tzkM8tFtyIgkaEnv2REvYPtL4b/wYdYMwJiKN1Eg/H7rG
56ibssqk8glkMeYSjkVeHp2eUe1vL5fyygvloAMgeSAkIWaa95G5i8mekLkk5XpSWWVglX1/p3pF
PxWZNQTrLuvoPQwVBfE6yQW3dNeuwE3K7DZfwo4fiHKQTRit1vafvBEsPWIp0XRbuQsWDEsX8x/X
dGry/zPSdZgp6xLx27irkczSVil0W85gMZHeAu5TVh1iVtHE4mhQ4NodLsRIQamh4ZVFNlMpF2qQ
qOoEnPFxzGZ7CRz3Lg1uxjxiC/De5WO2VgZol7hi+Wr0gBU3tWZAN/Op35DA400u+DWneKN5cQ2f
FLmN+BCmVjc7kAzJsWb+b1j0oMgUxxjSBVelFN7zfJ/WTOUTvYbd8drg0wfP43H5VI0+r00BtGdc
OCmSBRINbLFQilNvqnJAOtLSKnpv9veD4+nmI3e9AYzNU/K57M1bRsJXNlNf+TOFWUIP2JlRhJRn
6qB8dD6Db7Hj0AF6Jbrp6Sy2Kpq+TH2jexXaeLESU8Hm4n07Q1Rbj7jPJ41/t17jTrQjwd4lzTsE
v5yOhhCFcOeP5EvJbT5dwKOR1DC4CqsDcg+edZ3zqusPGA+Jgiz/X3m50JJTRzd1pLW0gfW3npam
D8gr/6gdKtdNq4aIg3zpFw4QHGipDs+lLaWFOfx/x452voPSfvdaLoseg2k8kq7haWoq73+N43ge
M1+xi6wHOXq6YBIjYI9wyWdetR4rY+vDoltjDzDlLHtiAK+wm1m8pCmhKap1vpkO401Jb5vlxqd5
K4JNW1Lanj3+B1oeD16FNKfVyj2u1B3vO3Nk0daiXCVCVofvxGkpVhGPanYVuHK8xZmWqSseoKj/
wk+yH2uXhigLBQr0wh6Y1fZy0B2lJPFLfgEczi2kOVe6aQ3SdynysairEPmRXosSbvhXpknO9Q2i
BfhIi/VmZDpUVuPSoUAuUBq96pT+W9oKgKMCCexwhgZ3vgiGw7l9PVbpG/Z01cVzrm6/n9SYVmiO
gn0wKb1gS+TGM/poA4/2T6QUeXK1xpRWAP4p0otFs0OUX77mcQHsIUeK9EMxYrF0g0b9SjMgmiug
/J/xh128NrKBTTGA/7hk1iCwaNIggfA+qRx2P0X3rtjIHlzeFpcKfQ/kTt38i2YIZGh4Ug3z3kG3
eHC8DQGBXTWj/PJJihqHOFlAaAjP58nnC6RW/EXNTUoJP/OckAliAf+5h1H7omX1/XMlsuPedcWa
9DnGq0Kzo6SXtx7KYzl7T432IxjZ1rtSrGFQHqvSa3dQ0sEA/febEuT5MvRtityQvGl3G/KDQh7L
NLbBXpgw+La3UEhMnvfr1YPYLQYGi18Rmta9Fkylkr5mLP0uRfDAzWMKV2sCaovBT3ggf0VbKnUQ
9yiNjg5EiMWhURUpmbOLovxSYzX0JgKWaBu3tmVlNnhFY4r6ZonzPSKn8ZYCD3CO5bFu3AE4Ux8s
z2xqEDFYAxZalMVa1qn03STi8MiNHPl5kaLcxuwsm0UM1qvppyS6kd5nTcN9bnXE/OGKlvAcD9b+
Ri7ZHffGm1IjKEXtgB9GLXgLxjrLA/u6s6SQVhDs2MEG5tPY2O8K6zuQP663ukGCycBXacly98uP
cAMz5jZg78EcFOAlV2CORHpkV7gHceEsMlmlBta8X/aj9MHRBmfBmjVGqh5rS1wUMNu8dXW6/yTb
Q2pca3TdlraOEtCi6BjplbQxsOGJ315px9zFmZJjJSI7zbVMGuwK+cc6LQTjg/5YnAtxmqiImkqB
jtfEsKFpNp8Rb7DmbOx0bID2ibWYYPreoERjxXovRmeQug55x80L/DV4iCIiJRxMop1aWI4MuCUF
sx1tuo3TmzM3CQcyW0tFKvMfJbq4ySpVInFtohstsRLPpUKGFPbowyJPSKhbp1VboHudGo6C0Z2f
9MgZ8d9xcuYE4UBIYAWVWf0w1wqLAlNm58AsXiPDPckR0jisgYYTY+nVe4edUKf7FHFc80DQyRs+
f/vmpSFN6OFxLdBO6T7HpeZlgV6zni/weIMQoh8zBt13XqOwvX2+Hjye7fQb6Jgh3IvxeugKT6+x
7mfB6HJHxnF2dDx/9HttcrVugazDViPVWhFdKuCrz8EjVNVDj2Xlb+rwpVXtHhJQpXJVAYc+cj3r
DrZACTm02Rm+eghlFkQieY9Xa9F3XaCenMwK42wdZ2E8UyQU0wFNAL97gPY2ylziRKn1lCgi2OsH
Qa9ywYWwyTZ+Jh5lNT3fwesXaLJnbNyPLlS9214BXiwpM+Old9WER/V4jxJ9WY9MpzcDkSnogHxm
7yX7y7py2bob7R+kAr9SlZ8OlIePPpTRvnP5GVekm6oxsiNCbLMkH2/onwbVSfbCx7X2jmMHrgD/
MEWoG48AoFMU3huPtKj2TL+KlshvmaYGB6LyttlnU8IJeQf7cTy8Kohe9jUU1+szr1r4OP7pOQdb
1R/9FiBB5DfoZbiCrXcOZEb7AI6GnWXDXTG2xuGM4T7TisfUJM7Y8xiNChQkFtucopATGFPmDl+X
myruNjItCcPaUVIXDBWQQeipkV8wvaXU2fe2EuHD25c+CshkHmaIOgNBom+gM1/S+e/rQZE7JPY9
6PgWSu0lDabJGT2hcUQxi2QKruG8TDK+YIt9+DQvJUPOBagzzlJGuIoau0RaTlHxybfdbYT16tY9
PfoxpNGBtrlBSXph20LM5Smt8HNlvsg5OdC/mBZilRy26EAjSeFDGlqg60Qqqqk1XMaNphimXgLC
v20P5TzqGzzG6Ma8tXnRGnIiDRCQRSfOlYV9xs5HwJmgIWb+TVJbm1p5IfM6WpXZmq1KMg6i7Jy7
0IiJfjwOpydmW0Rc30ghg5qJ7h0i7jXBSL0NlLpzunQ96SMo99lDpgFCuOromSfUe+R2pFP3J5a7
xhMm2eibkJMozlkbOhWU1avK7TgPH1b7nixNyGQmoUqP9VRoDYVgc0C01djGeUAj2j1zKk2zp75P
Do7O2ylCR45HSRhQKiLVWMBcFk64ChTfTN87nE9jYBTsdlBe4YZchB9NP6n9wFYcqUhUqtNZL8u8
gUZLuw79pZbv3oDdIdQ877QZtj+wetRQxiE3RdEcTlRGiRX6U2RITRK46sCscUO54kiX/F5r61+j
FXReloz6iGSHcRl3vDSU4ClksmF/avEGcb1JVdZxjPnPSvkUP3LHSW5VfM9h+L3G0pNRUcvM+JxY
S6/yqNDPvZId/Iu2TXQHzyEy3HrefphcpLEiLXtW1y7tsMdvcPqMH1R0Hck/WxnMhatFu6gemjwH
FLrnCHi271+DwhU1Fl4K68g0o7EUzRXmxVYYLFBXnR9WWvW65dlhsC2uB/s6ug9ySBJ7a+S/cD2t
ihZgnsaI2VbProJ47awQD9WB2Im3hg7OfflRbYQheDC6hZYpgv3qwQcU1+Y9wrjb7tDVWRJ1xsYb
mSUnievY4qG+mWGlHAWbe3EdtvDzRyyFcDJVxEbECBlnsmdwMtKDQdEQ6hofBrqr3YvmNoxxW9Qy
cTqGPpECF6sMyKMlCzXNh/uPxg9qoNLmbogV5Spk5/fWe3F5xWKsq7rGAsy9GZeAdo9ls1Te8/PP
dvp9vHPphESOA+TL4che7nVVIcvWNU6nTp4ciVMWxthFVi9YBMcCdjLddf9mBt+oELH4oe7Xj+ub
IVKk03kMPnlGvru57hL7C7O3NdqA4Jl8oQdZY/znAcLpsxwz/TBXW4uG56HulnbyQixXmochWOIY
DTisnV5qu747LdEov8CASqcmWUERv+KrafFSy/KqvMOzuLWFnQhaeUlO8pa+XiiKeefv5PjTBdph
a+OoXerJAdIxmkfbRQNenf/7T+H2z4Ywf4dZSUTs0LsRyuqOWvW/MEY55jw+VWeWEQrOrjPdpqwh
Rs99Jug2BTHj2bzus9dkB5CwASYtNz7SxbST4P96I4LMbGxgKtP4AIQOyqprqVL+3mMz5lK6+hj1
CDzPhstlTQwuIbBcaM1F/l+OHV2TeTZ+oD9QpEzU5/OdWSHBPtkABDUct3Uu4ZIBQreUihZvNvtv
g/WsE00I5kBCwMhEZlG4fDBcLtEriHz/iirtw+uh6hx3p6xw9EhVHB8pps/sGlwlT1uMPMCyIhay
JaQ04Q8ud8qjoizSxUpVXegn09lvtZh/3piFK3v7fVfpTPMkzhVAmUUbD21EiGEd7p/rvEEZkD+W
VFXE15WY1zWnf5GIrAWNh3QNRZTeyfGaqOKEynPu2NWVf6TgR9+onU3rQd1xYZxcY7Hk7IOxnpYs
NJFqgdlj5YhwGyb4/DMj8I2Wxgc4e0bGgPiqmYgiZZgl+wPEjuvhliWm4qXx1WsYm03+bYb7rn1S
u9tmCNt51R+tNjoG7gBXcmmGIxc+879rClavvKX59ZGxJXP/Xgdstsi3B/oK1cbCenpuO32IWtXA
LyJw4rhuHlwU5fLhsePbFNnBCzRQvaB4N6XdPh0DtfYxOpfl1ruOt+wLiLZORg/634Jg0cNjHQkv
ZwXiRmgotof1MPjiU9hwnR0z68ZrOfkdYcOrQxhyB5zwMauSt6TMhHhNUfV4ewT4MxJmFKqAevRz
Sz3Y6at0c9mwgDSHBMb3gec9zMzFeXbO4XQBiIXM6D9UJYItL6/1E7iobTDKthsIGx4GdHQ41VSQ
yPbN08eQzm7Y7VxUAkdcBYOq1kkkzpBewvpCdHnO3EiIyQFQK0dO9qHm+CYcLWxeUb8hP4F6gdFW
h+22akEJ4HDigptUNXG0Lo60XViYT8D51ROCscKsCyrvvOm5I+y8Pif95Msp8O52udmnYdhT6fy1
/9RGYE8DD4ABEhzecdWaIIDxxhVqbDQhWE98g9UnBRNlk/HHNbLZLy+Fccm7UAHbg9Fr9+YTKCSD
qBE7Wcq2v9Vxvk3cl8ijGHZ3s4JTLkG/lRYcnSvHOkedtGTEUrsnEDzzSbFHyhNyUhMrng2Z9tXV
aRHEHi7LQhx+aLnKkwUoqe4l1UKRbLhpiCTIn5p3emeMGPzLbe3IrflMOQjXuHfOOBktz1BV9RJq
qOZjaQTFPSvGoqAIKlNfp4RPWIKHBspPL6If3pcG7dNgo6rIYd5xVT+tB43yNPikaIZSfFQZz+UG
58hP49dVpPObCj5QKVGUzXFtrFoYCdjiRjBPkuo6VBDkvJeNEeGX0RwclZLqHr3JeZFpjb2ylA9q
s4Hzy3/27Q0IXRZG0lh3vNXJ1zsAACt7uOsYLr8PDLDoPQnQ4iuhTz39uyxQR8Pwhj+d1EY3dotI
1cMzkkmLmLWajnNf8LTYKwiWy5N8pTI8OmUioptOzFvEKwJWQklJxR5lMXy0jcnJp+MlOJmW5Rrb
40haZJVLM5X/Bobe8+Lo5peTzOlOOl6cjPeVeOeHANFkU0l1mufW0ngSG25tB3ALhJL8a7ZjaT8K
9sxWoc3o9uu4BPWuoND3m/aF9MP6Igkv27a2i9vpTwsUy0X9YNqdDQO1ScRhdcCB00sWW5IlXDQ+
8oA/VVm3LgwNi9/3MeoN14dJoi2xgZBB6wR2DY2F+e3U2awfdHhGsHsNtk9UlQvCjLubJmVC2rkI
ahwmeGmXntcPBMdWFufGeUiLf/vgjBd+qFtJz9aS8+6WXjUDR2oi+sT90gpiBL9F23yIdAcSv1Gd
mmDVPvtuGnlrNB+47AWTyl3z+eMHSp42NisHCGFzv2B+jwweU8BIM0KytoPy7JBoNzmJTA7yQOMs
bGuRPm0z6zRHtgudHLPkSw/FZzpPJGnq8Z6wNyCCafHABsh5mUBpPSyOS6lwVQYx/aTHYpqnyY6U
Mo8yUIsWscx4fZkXi8ZAgTl4tTVpchiSYYq+GynCqDYyReFc2v8g3MfwoPYvqkDskIC5EyPK420s
3von1kj+rA7LkqoMUYOZte7/6qKoJzN3kvMlbPmxcmNN7NIPgZLq+8h+2beET9j1HL85SufDezdc
AejeNFJUAqgUlOCe87dggRDq/T1OjxvgFQrYqIPcjtnWoJPgpdlRvtb7OTz5nXk5pQ1DRyUteeMa
+0672XOmyuHQXcZ1dEB2Ps1qVk06Zg0Bu2VoYvOXeHu97VTk5VSzeEVXha7VX7v+LqZ7RN36GewE
AiC1bzJO6uP1zkLWoNuOPgTL/Iw6A3+uEMgCT78eWPAJwjfaG28A32hai9jB6aiRPqEccDTuWgc7
4f756aRk99H0H6qOU22t7QWtGJ+fnxB7RKLtPfWaVhKQPpycRd8D7XMT70AyOyCBDkvYDRFJt0r7
OOCKoz+J8AKN+E9ex0BfIINPl03crY+nAML1VH7TI2rioQ/Lxd2rkUBZpJ2qOgOAcapJRxjLFhu9
mE8dvWsJ/f9m1HaMdw/cVKonrhVIaBsyiUeEO/vJFI2qqx+XqchWe8Tsbz+s62IIVl0CLpfC4oS5
XHmIfsYsPfglOV6n3TrYfC8/f5ui/OgiV7sqQBdiYuUbFB5OCBNNBZQZJzq4KMu8weenuHH029+Z
EVVmqYbkXVWQ3lGi0J9neGhhJQ0HL38ZyjxdYC1DTGrA0euNVPp8VDSoZ9YEEGtdfKXaNDUADRwq
igsF8b5oU/sqSBZEDOKYfp1ZNq4YWzFxZOY+zcjEMWT9pL9fsJ0mYwxgQkAyzpZZ+k8G8jIkbE2R
ZAVY5r+HiT1EVEbl1HFCLZvJ9vygICf+9sX43MclSHddfSjVZtKUt8++BXGooNi08mlgGPb/fcyV
sjoES8E/UrWUNs/tlbdpx3anC0PuGN97iE5apHwinXguWPRRXWoagNCsh4pnD6Fp5bG7r3MiHERG
fwiViYqac6TcvQsY/so7nAD0QpjGY9RAZGJbAKuCKnqaA2RoWgr3ofC+LKHti0CJAy3IgPz8rwBm
gYoWKerfylHulZ9kDlcKcanm/E1LgWAMorHMCZItKgldMFWBeu9jnwbnVtqHn1Yp44DjSbU3tfxz
D4zmQqE0Fr+l1wJtUVYL++wb0+gF5X7QOWCaatYBBWqIMTJDJQFvmw6kUNv0t9WM4Do1gwNGXx6c
U6jzIfpbMfAaogtqS7GARS50TKNPIwUZnYEp5KoEhffBSlnEUqzsTQW+9dt23qnK3Vy8Ow9VptzZ
TshXPrZmyvgsv1b264yRlIpxNxIxQUFSZDV2VCdOuJGGWWr0iYHOZCGTxEPBsL2BqOcOR+yqVA6W
LpjcPuEhIdXY3NRTlzAIkddxx3aPTQw11lRtcLcH7UQK8mMK9K9ap3nvHBVek9btyxCxVwwDwv9Q
q8J+vXdCuxZGqLXhohwCkIn5/kN1XJRk1bZ8EZHDrNA/6ct6Xm3vmE6MFjG7PckM0XrW+TcrHNle
y33Y94Ij0ALDNvVFMQQXMG63Pd5YMvmno0/M80boNPLxR89Q/6V2ymG5WZY6OIUE9klo67KRWc6P
8FzyUsxudetkZDDF8SC4qNWDbjWmCl+FVXXdL402p140JQerjo/CqWbXY7fN5mpnsr0KGGEsveR6
Ta56I6Pt38udF47y8XL7urutc0etBPkZHlZrcpotzklGDI0/tclG/HVTECRZ9WBejFxpITWP48Jt
5J72dRsIg1LCqowq6a2DvFicRaXRKtu8YsiIQeGtbQBRes8MVDSGN8X2HXrqleDhEkLs/1akhPGN
EKA1oEjpjP2zYWGrsyATtVK2N+fC7/rwk/toDbsV2b3J/Rt+yla7UL6o4+OcIjwVCgLCd+Wsews1
thDVSmdKgW5cBYBmnxsxmQQbvDIAfRN0UboGSv4FNFf+jb52kGlT8kLK45w0HDNEt7YFjjt0ZsN3
UvYcXutt3kR9uFbeslCz5sC/PlN9+Hr+6hNUOgiY4tORKXzFgXNZxrhsIfN8byVm3IkssuFDqCyD
q4oOjh6ljb9SxOHpYS9JfIs5Lp7XNjctsh2GZQa9cJpFL5myX+usOBZBhtL2YbOAoSKBcN70uTBH
UEkE8595x5gSvUNXzlZECEOctJ3L2xjbcHDO7215P7AVqNN0ViBX+jWs39Hf8tKFJk2v4Y0prPew
OUPx/1bP9GSo88GRIDm4cEaFAJBzmEidO4AKy42zLbtLpdIoBA4XwcsqDiIrtx39LUiAJ1L07vqc
JeJPPS9G58hdABqhJJecMirzOInz2EFI6d7HsiFrgrIrKBLx+Il1M0Q8YOvMHr7heuD+igaodmUU
0znrbvTCEH/Pplo0Yf8ccSyHqO9I2eNwf8BBNRdzgQN42j3GKra7yR7UUC7TZavvpDJj9cI2kLS9
5QVF8xnRSiDIVxRkt3SuRbeeHPZUb3MBKwSB660XPyvxjbLGolytOLiiSdy2kJxQeIscCGgm4kvL
AF3IAPjurkiLhnbEo6+own79m2Idg9G8ImTkBmFJMvj9Kr/HU9o8JQ0KnChCO3aF26fY0zVZ6tte
7zrpAuR8g9Sz+ZNTlPFOLvzHhFwwHVfrBjHxo4WKY8QSWpZqoCbSMGW805Lo8RBcOboasO0Fj9mA
Dh73Kri21zU2WdPoFAFuLN8MvW8uYuDsJtR2zYaclizDEEoK11wjgarc5zlzT9UyPnUhUDqRU0Pj
MUcizxwpwZNO+wmX/hDdBAbS1gXAgcIfd5TkRM08UJ4z4IPm2WhTnDHipRFHNnOl7hlijUa3EILR
JZdwQySPmapgTzG4vPjxtC56dqqm+kwaJfO7VbMCKwI2RLLSyVBf4x9yG2FNo4R76braucnaGG1v
owt1hscXUHBck2BJoaHfNDetvRlliIMUveERQin7D65895hiOqNSXZGdJD5yveHMjyF1U2MTmyw3
c5q2wpYPF3q09JZIYedqUAm3nxSe23KNXLS8gZoYjvreY1IFfJn7AccZnFW4pzj58qtXSRtgxZC5
peAzE56ZWpnWqyrN9+q+12GM/Kr8ZXWASfO+/vgIH1LwBH1qxq2zXzlz2rFKaWd8UeqIBvC2J7O3
4+MuTINNHfD4hF4H5Lo8boMsb72K492/SoTVAXjBtAqfxUFzPKjSSDLsyu9l0KbGnZRHu7pbrNdm
85XtBegDiY5E9U4628aM8sJuZRshRJbB7iZh9SC7TeV/dYiAu03gQi87pxFXP0g5WaUu4gewcFbp
e4Bg4EP3qxkD9nmDvkCdkDYnJHp73BNQDGFdnLYdtRiGuJ7Q4YFU1prX8tZGF9e7qw012NNDe1/7
ZPkbvt/gGeuPXS8f1v1NCuGx4aXWpbjES4rH4IehQx1n2N61XACwAa2A9FQv161axJBOnu4zOlCs
f6dTCVYfSHJuUgqB92O/q1hGYQIsptKcxPKwfBdYgVlj5e/zMeulZtJvWTNY0ONv8rgDa863VKf3
fFsUx4ACdGOxbbMWNWLaBC6gDSXAnnKXnAByJWA1gWZgMGeCxx/PMnf/VrgL2p7sleacoxzBhl3o
JAMrB7VmBT0cZmUeE3E9HPqjODWWuW6hlIrMn8yElR0kq0Ue+7fXbAdVQkSYuCLKWdQbLrRER0au
RiBKOeGT/NbSEZX1qcQdGxzoMWixpi+X0KX614R7Y0GCr9lVXGjsIufXoOS7Nco8hfxJQmvjDG3h
08fNm+W59UsPBRUhf3xycEAWXSAEyuONg+POMPOLD/ojEfb1FlD8dvnkJ/VxdwG0fix1w+uxj17w
ilTRHEUBc528F3cqGeMsZwCx0jtGUV+IsJQPBEyEbT+atIv1pOZDfIMcHr3zZJB0UwwQ3ZngcD6g
EXkSt0S8MptwQVDn7KgiNB51mTXUb6S/1HvPiYAeY9s1415clkdD9/K733v8Leip9kVAwpshh4Nb
qszpbtL7yntaeOJS6PYBe0jDgG/Q5lxus+RVTg/33zOlfKHQ6gFmRt0STS55r3rh4/nXI13B+bH2
azsNmjgNrnjvOS+Kj9EtXKVjPAx0Hwmt7lfLAm1d1RZE1bHsawBo7+y4zx+41w5fozh8jb+RIGvi
3cpIxgtX+pJn92IuldM5kVEWKc2QMvWI2h+pGjavSflSH6wPnrRMlFcmQQ5kbdjDJGiG3G8QF7vW
r0BdZF7FLMeII9zDpVZAXKDpsW5A/Jy8z/DElk5VyPxsLKR7R1XisfSB6DQqYXy2PKQMU2icpoBt
dK0Klf7qUEjqGcJFy09PV6LWpajL5+xHSDwAoxwuT1bRpb2ERac1DZzwH9S2yBA9A05MK+GBx35r
/3JUqrTae7j3S8Y1BqJPumEREc2lUGI1KdwuswEFnkshQCzlQGkDEMrxnHf6P7A4dbib30SAwkAV
yFMxTn8YZe/QLZLxZXWe1k0urc678gX+cIm5GiqCrkcbPIIunmQjICBgKAK5uKF32rP09o3WZ8uG
pZ9D78K1tNv3MYjMPXFo7hH2nKnWIC+bC7Vpi6tIvLygFmm1RB6XjjnSFnIEDj4pGksikw2qSLEw
5m2DbreXIMuNDa/H8/600Xm3QsNLVkuV5iWT95hwRibzy9YAsKGbOpV2bpyBRFJ47gvTJhU4EUk7
TslMKkGZcKB8EDaL7QnusArC+mHk+0SuJ2CjALUQGeBon9J9PppVd7EjHDHpSqjBrCwSA5eYjl7C
9sMMpZnTDDi0WO67sZe4LfNtMAT+cXqIps/s0FQ/+HfqFhIz1XST1BMot3Cxt/TRHeQz0hmCqC28
XVPMAXg2NaCN7sSzWHJNAlvw6TuhhGExxV9U1BHgrpt5AfHDwlOFRQJinAcb9SuDJ0cXAbKikFGC
VR7oOC1gM+unjg+bpzNomwKP8WzKH5XMh+1Vqj1bFzyZaGcuQ2mMoWOlV9hSsjcUAZ3xzoZPVjJ+
nGU6Bx6qahxarXqJSbdaDZa29/y9IQb3L5TnnUPJZ1xe6UFjJ8esUEzsHxSYaTiFz2bAo8OhbYrV
uhkwhZZN5mlLXHebfAY4+3E/8PgvLqntz5KyrOubkKQOvGrIz7TQQk2gO4VpTivC8z/lv3dipiBG
WfAP/W9q21fTsMEdniSiixg6wZPeNrPc15YXrAAPe56KUbrHbxllx8xeK+ZSBnzrJQKiROTM3OOO
gCCKS4fAEMzOjPJ32JIZvB40w1DPT6CcyyqkED55wFHuTYesBzS/za73BzsCX9kOn9m9f6knrf6O
aq1w6WvgtAEo9/UVTRtt5PWKD70qD1D4UXPOWtbtKmML/VIAg2K/QujIqHhoJzL4Xi7z9cyTN+RT
Djj04dqwNerKEzfMfOEtyjTFl1r7fXz44KxU2GQPj6CJbauq8aywfoE6uJJe4A/5NEzdIkUQ2Hnb
/HJXZ17psKM43DfSGOfVwWuCjQj+BtrXlpEA3q3ZKxHGGRNMofM4Pb6PZ0AT0GPYCFIP3TIS3RyH
/4YLbKbmHW2b7yOS3DzxW9cNQlWyFHdWz1y4JKR0keS24NMzR+oK4C5MvafEpAXeVp6GkuJUxXql
XQwdpTjzhXhMHShl9j+Bz9tJPSqn1jwPJhJTSfdFFgz+NnLm4MGC7wc2mFnqQVNZZoxR/e4kUPxz
fQA3HaFWPy5HHPkEUb7nSzqE7P83t2DMdsto/BhHquDHegdnBDADf67/F82DCnQZwyC4p6jIF36f
2MxFdsFkwfi9ZT/z8Nt9r0ppPuJGYdRi02ThIVc2hI+Fd+I3I4sNf0f5j2n2nPD0ZwOuZG+QyLbs
LMXur5VTJFWRDij1T4ZCgR83OTexeswIGO3g2oGOIZSduoGLuXTc+oNJyagcT7aHKRD/bPvve0AG
QGR/KXOa0gn80ji0OXZd+bfxq3asuMTKwPaWSOM3+uTpRrcOVVaO0oh4RzMCmDP1pD2088thnuw0
C0Cl+lhkwwmh8LcUUSh/6eLzGMG4w+G0lc50EUIgruQbtVnl2JPw+pQMq6TQfe85MwyIiFn4sSqT
6sxn6IURjoA/O0Ccatv+d+0L0AwoWIy9ktDLcGAfucxbuvL0kfrcATmBvTEhFwotdbJ/VRjQ0OQI
pPYp2vG4kBZQzbcIoTT/fi+KR2yOOB3BS12SoAQ+CO8ayJXjzma1tQQlk9eKgXmae1io60F+j8zv
hKSCy3b2zD1lZ7Zux/tU5UjrikIJGWT2Yq2FLhrDBl0yp7Mzm+SqZ4UMfJVv0MH1YJIke/ylMxwK
QaG0BHWCTbTK1YxGmwvzNOXGXehH1xrYDGkeFFx7mOQEr2Phkw7E47bBzgrGMmUtWsMfQ/GUVyxP
qFwzwdodSeMLei2E2cPLfIkYcMbPnbkFiopPNmvV7SpPRDZe1rGmZDiYL2wBnD3TwkezmEjEyLA9
Pqk6gI05LpwvYaqUb4/5tkhwKgqiT1oIXhAeMgtL8jYufA3+nU9776y5qf8xghTyfjwnerc5YgpW
+3EgxRwkPkkMjg0SZZr4QT+c8Qa7ungugwiYdLnSTCe4QxWTX//tHaAV6h/DT8mR8KsW3uYe3IBL
U+RWdBOdSwBZPz0MGIA0o8wYWLQwE5loiBssnX2LmZueo3nq6y5EPBBg2DrsU5B5x6LjO+jo/IqG
cZbujz6l9Zz6neefEy5I+ow9rIDXSyJv70GUlx8p2GD5JE8phAFwRSRcJRD+lY+4jvP4yyQQaWuB
NvuRRW2KZa30YAooBPCoM05QW/alroXzw7V6jt+M8nt8M9G8JLuTHpvvPvP5gAZ3jOFLK+8ovWKV
2az2dHqrOhPMAlwEUXSe3+o2/LT2K6gknlYemGB7+wloVEbGyAvdFdsbx5g9W19XETfAY50uQ37w
s26GW+cEk//Ir3adJfvJYQ/yJso77PMH3LQDvQkTQym3QbekhVN3RNgkgGqp+fwJvuZ9faJjvfia
3+GRmOoMGbQZICWjFphwOmxXmZPdGQSkwkIoD9IQpn/Gp+SuBWjGUM0jT71CZ2hP6N5oOf5Wi/AB
ljf2L9i4uEW3nQX/IeN5UY6rBhXR1k7Y8cG2U5Tc/nUc+5SiT0Dt+dCnY2eoQjVWV3au0fMrxIpt
upojPOluAFHt8JmhYCmhQhgxgaI4CTzzvM5OIWcLcUBfJIsbLOdRkQBqiF02KSTo+R+ip5afCOuw
3Y3PvUK7RgpsJJsperIUh3n0mye6bQ8OKTETR869H6TiW7p4bZptx6ozTmwYZOKCOEtUAkuescFf
G7Sn0uDvMCF78cqLpEBw/JtIt07t5fgDWn+5HkwIFKFo1ReHKHNJbi4X0wiErDIiJTCmxecSwZrC
Wg9AfyVsNi7hGLIlfldtL/ZebkpER9Lnb2h2ZbpBAOMf4Z3+9FdorrDoerwjqP7O+YvdTzNHswvy
pOSYrf45eDE28bnMU/EpZMlxVkDCxirXiHVSLNWGvB7g9yHH8Jtran5pO5byBR3cjnLA0On/n3Ux
TDq6WL6G9X/l/EZsTjFw8vOisFnlUl+tB5V9ZF5i/YXolH4fwpkW2cEPfZCa6s5DfIuHDkJ2M1DU
0PUxRXwacKK44iSIvmrlnpGDMaMFkcG2XXNDPOnT90FWMSJRV6fVsHulddnVN+gdkz7+oEG25deQ
DaHvhNvFDZP2jEGabhBzxfSHyEzXnGpkRnY5i/dcNLwLNrM+RVWIWrsszJ8TfOMuo5gnzekuF3gu
ISGwki3BFiFS8bUqf1X8R8DN5bT9AC0F4GHz6tindmMhLrhz+U3768Y+zchZ1OGi0epGSuYpIGi0
LJF9w7nGYGc50LeKWccasFzFRcbRIVE8oH3eP1WCDn9+BW4n8BDDv12Va5DyjRNoT1Kh4WqnJLN2
UHy1Y9BkB4IxbhtyIRcwAXXhoILrcd/HfERRPTFbfN/4/nAx2ppvjg2XVDwkrMunYIgc27QwOyzX
4Z/pT/+OjjLJGDULvaTdqYZJ52g+kicmh032GU0Y8QjEL4opfEv76vR1cpKoy6h8V3KyrMQyJBIw
SGb1bFCcaS0Zn+nReyAlLXrV7FZQNEhGCHiR5QtFhF3xUBfwL/94Db2o2U2zt51+P6YBJr8AQZ+K
7JM4w7GMI48oIQUMTebqbnzWkZe3dThY4qPZL2rs1KDPJqJBl8RY1ZCIg4My2/HLyVAAcWfCWW2M
AmFSrQSDogwbc7gkaqhExTB1yh3tyd6DDzpa+fwF9v0X6aIZzYoRD183/KnimOtd2Ci8eFtYC2Jg
iLPbac5LMUNMeswfsz7IeMy9ViuxaT/flQI215vAAYg2I0Ke+uASnA0RX4yBTQJLBz773mLsL9Up
mVNSC7P2JrqQ4cab6BqxLvhXwr22sqJY0FeVnuZ5Ux6duu314ZknmbKd4CdhZWN6CrTfVrK9c+6+
I9nlU1/bWXFm6yXkj5YjfNqrxtkmRmaOgYum57FFERj17z23RpoHGg/leAMAVQtdoyLB0OJzYJB+
a4mDYhCh8bdrP5RqFrTbNN7nHg7cZCxPD6g4YgFoAel4tPXU2jQTEG6QE7ICwMe8IWT1czsmzr4j
S+tQ550qrWcJwPpAA/K/VZKE/9EQuB1g+C2PTCtYPej5O2kt1OIIQIx54m48PhpAkeHYM7Cf3pzF
59Xbu2oDrTa4HqIc26SpY0KI59q0Nex14RnyRtDBGwYo7tKfBIe/13rKn3YuGvVf+oY7p/tZNtVe
7LL5/FZDEilb0sg2VD51I8rWKEe858TyhMaLIdMez4ElPLwj4zcf0E4i6opYZphhOPUDF99wbSi3
XMMFODkKJi0WMKRwFMfvf1M69iQodQyDcVcod3f5yVoCIJ+1cRdw63lkibrxrRuBG+i5VI+p2N3G
cadjLuogMvtsPPE72pRQQkftaHHwnExtOgfe9G5P9lRkWvt8PdxTKR9UYG+ztFUNu4JVuQ+wThhM
3Z+hhzbUWga3NKE0TX9ySTerALGc8Az8BTMzk2rLrUC7jMzvalE6F7avGU2q04X2j4Q1I/NLpe0l
NUgdhn6ld73oMRTVFXMIRtYc10AtgZUiRZyHbgb12MFTOwDntBogASLibdd1/6KeNvKSYCX4pKgq
04G2m/MAHTSwFeRwpSdZXwccM/41YHpsra2HqjawqFFGIUX4swjmGRhMJcCZ+lwDsz9ByOpFkujD
MJafzWzXP5p2af+sPDXS1bFGhgB1pbg3EsQ+MXp9oC5fbXYfDGBe92y5xx8r7j5fp2/Wh5bWWtrb
GqX1kIqBWowp5gnjRehBuPgr14NMhTGmLPfGy40Qw8D2p08OscCMoecN500zRI2vsv+mJutjo328
igNhLl2L1Do160Aqsf65pV4bUWHiMQ1rwC6rQDbHZiGU82ayR3/n3gzssCtF2Y3kk1oOtSWowgFj
6U3ZnjvXffphyfN1lG6H7A8WQ6iUeNYPYrYxIbBeAVlVX/3evVmZJEh17JsA4Dr08qJZhzmang/n
l4+JTDMovdrK8zUbFdtXdx8tO1wQbL+WmRwcROwxuEWbtLWZzRF4XtbOPbaezBWoNSuIQc8Z+gPG
Zili3PteoZ+5sA3Iwad67pNpMwpHL23s35fO/KNlEHIvBQFgxPGI+rdWy79TtDxwgpTisw/+DruW
UbH0m6L62y2gg0qHdYJgPPZLQMo4HuTpFA/uPb7V7dtpGeUq4SnV6Fu9zysaj+mM1S4YYILgI5lP
4gj0EZrOOKsatDDTu5jl6bV2xyh4jkwPvbVn8EeClw1eFWQ68ZCkI9bkAOGVysPKZ6gRM7P9UV6g
1odb/WASrLyQ3I9260ofebTqWjBUDzK6+vLA33u1zcWhrcjdH2w5/YESzpuYwPv+bnHQquPF0jpf
q3x0vxqkR5eXEjkNtL19NWaM6BMZ37p6wI9CyEZfW4Jn6gW1ftqrgr9VdkZwyTzkJZDeP5aX+1FH
hVAHz3a42BYpBOqrRgCj5qHULUsZsSfaasVpcHgRQJSvCmL4/a1GwNg6cUw02+tPLiEklb+bNo/g
+mEnTcPck8y32Zva04AGHHOrKKJIWuvciD24d/3aOffkg1WgVOvVgF/EfHZjM2rNtdbBjIbIIRMC
Fa38/g9suctz6F50w4996VyB2MZSXfYxt01H61aoQfiyD01bPsJUSykHHFRvBhgWCV31JjnTF40a
qFMlVk/mPUi8aSEU6felsqiaxLjeY0MfbavPa9AYpp9KeWEMGHTw1XgqP0ipmhuDKnLRydBO3l9a
m2mlKYywQO3jd5YSG0APfbg8PkQKaUCg7b/xRv/UXjWce6XE/ymhMsERpYE4Ug0t5r2CNv7fpdgK
HnvH7ah9uxZom+8cxQImr06mTFtFWsnfEmo+0TuL3FSAYOk91mQleou9WHHI0J4bjrfN0lYhW3sK
mmdsarHZiSemehXhp+6GKh3e+8DXgE9aHFdBoJyAeu9cv+UkLlX76p6oKcNHG4Nw/DnX4aTF3nxF
f3uikgex9BQiznDj7A0GucPeXs0RKgsfQQvGmdR3kdP/Ss9BPkNsO51QddRtnEkZQWYeMzz3DqMe
Lq83XLroBizYJgy0p0/Kmq1XyjlDxNd/fyx2RyccR/n06XweLZhsq9liTqLQ3RJBe63ZKBeWN9kD
a9Cxcxi3O9FYa/8BgCwuTIsbAPgurQ4OQGVYYkIgEUKfulgXDG9LL/R8xCWA/MxNcozc4ec7/FQ8
mX/RrycpLNQQTKTAXmnVSnfZ3zt1DGcSt/tlYAqjTvVQycEJyThIGJC0NGnwSzdwbNBZFGJNwoXO
uXN+GhhcLIVG52fN+Ir+sw/QQshHpMkbT2X/LNkXDm47spZh0xfE2NUeSiBXZlQWx8/CSqTwKlUZ
HInSffm7/s3BO2uTFoBeCyQ2Ab+wu4gomdzhAL11tn3Fmz8Rg4fldfH1JHsQFSVxo9X63FUDVKlg
IugZRfI+CqmxeLorYq2AASivsj72Bari5S02U0RqTLcsKbLx6cpN5XvkZV50aHgbKRL8oVFEyAS0
shmPT2h5mRi76xrnhMiccAtVJ7V7Yjr8uxzqrN1men5Ml5DfgUHcqmkpqdpjrQtnLMHD/4aJVUCu
qDGwBfpsI6lx8ArmVNJQPut9Y8awefLwPJL+cqELaftJknPJdeUO7JQAYwa8g3R2ml6zCkYK0tuf
IUqNT9EPXOYMOp5plTK8QUchZ5xaDpb1ZyR4GqTrCuTmGGZyzqT7F6kTfjD5NFwcndVII/iP6fOy
Ljj0V4mxITl8dpFGulZD8QtWpJFLs2r7LUWfSgFiIREqtC1G/Y84vcRCIwCiKF64maAJRZadvS9X
f/aMWbAuZe5LIruE7hCzwSr1FHpqP1hPN94igbrRdceIAsRx6eKqLVdXiCTYRySg9HPlx1yCFoV9
6yFb3Ui2ValC2nziUmmp4ZrQEdioSXNQj6Vt7dTyXiot85Q7A7kMshteqj2F52uoinVI7IVN5rA1
tz+11FyCoNDbbPZj6OZFjIKw+NcWIS2IGoOjINP09NEnt7BFAVwqocbHoPbDPUbiHopwo47aGzxJ
5GNysgsAj92kmi4BaWcgM/pyKL3Qlqhvc+zjXeMFlr4HeTORsofM2k2HfaVtIgEOtrzX7vGopA9+
SOcGY+tCU186h/wOoB+vme2Yo+fsc+mltFCYsaE3Ee5L4RLR0JTNIJLzP9pXPNGDPOZVZ8P6m09S
X6B4A+jnTZvdcyX+wZZLKkYEN52o+IlOb10msjrQr69cz2gZ5566vfn6bS6AT79FBZjSgSig6nk9
nEhOdsQlECoh/Uh2/4z67m6ZYKERAKt0BlydrNKivymWcdKGFTUlLXxQzg21gj4Z0lzzkKAzeHTV
jOvd7FWGpjRfV41AlnTI36mp/AYn0GudTJsm4Dox7ES5uXouhJT1tMy1e6JKzx8JjTgu6xI2Wxa1
iIZpbySccYBgjeOZpXusCGtQjA3vaLy3qWynA86hVNlrKm6odyA+6no4BMidwKNfouw0Qo8KNI8D
xBFkc5ZLRccQJpqe7UDmQdByntTcEMfcK+ks4RbdEri73ARXJ9PFXGG71y35bstUOjY8Z1gSpmFy
Guq3Hd1hSNmtDOo7Bb4CgNDbDXxubNh8vAtn9ke+4kN2PiX+06P6564P/aeKF302TFdpHbP1UvV8
IWH1ENVbQDmaf4jALsQ3fNFCj1rAiURo0dnPQBk7sxAEjkzyZMZpAUvS3kosoniuwrFlCAd2gMpX
dhFxlDqXdIWIoH5/Gnjj8L8PqKF186ymceuaD5E0M6GLQR1xfHUQ2mSiaWGxAyTyOiXFNlj74q7S
UmvQmqmYQ4Bjmhmo3NFdaDQMb7KqyFGsn258+klpGj20EW+zb01Vm0zQ3qEDvdIfmFsicqtQS83s
FPu3aV/RkuETfmiWdpT2s9t0s+NQx/oPxu9WwivFNUU/Wy11Y0lZHaHncA21JEqPQHIFsfUtG1D2
8YXGwLjQJhS6hlsC5SB1ZJH0CY4ncCdK/JFg9yNm1nKDJ6W+tYKwMRe7AE4frdQEOfb7pvahHhrs
hcVqE2nKvWlv2FN5dNSRo8l/ipAX85nhDwph2waSq7WoJNVd2neJzquOf0a58lXe3yqCpYXn3euG
Y/blsJLXxlqRu0g64X6X9vf3pxymRl0RNzxaFdDC0GS5kV7Lv8eCFvzAFGqp5NTMTbd3lmhFZXjp
M6f6ImdS95cFeuJ2p4jIGdkDyg0lNVPbuEX12FbW5fvNAjImJXU+ZurKeOq4AAHDuDx2qnUYbSbM
h+OujIM0bwaPqGf1gWtkLKWFw1J+Cj2r8VKHwSI7FaOutilbqJjpj9eh2joKHgvdpWGHc7LPoEZn
RshlEZkiv1noe3QuxFeZjDOMI7Vr3IiQVh/HaVxTymJXHoCtVSWucHkn0uWxi0QxMx92gbMeAq67
zzourTKHZAcAser1Ll0cM8hzh8+kmnCEjf0jsl252Ni7BvE7QArI94bhaKpgtxVRQrZ/foF0v0WR
z1rES5j/7bCQooSpa5N63ob4LS5iVM3qxaEgi7Hr0WqDV9OTIH42K8Moq867r+7K5lKChf2trkx2
EN3ZK1fFkza3I39jPO8F960l3wo2F+3TbEYmsme7hkqgHno4REM1MH3/epF8vkDGRMHO3DR/xKdm
FVeink31S6fm7JBxHX91WWCVgec1Gm41Fm7nSlkrQswOo9jluip60HPbR8+Qz4Qj4gKa0EHnyWNy
e+BpW+3AnBKdhNPjGQI0zg4m+EXCL0EYtZtLzNBSP0J5bJgQX9RoYzVPiantNnkrfiAEO1IeRv06
AnMKR4uH7BHVhFz6I9wS3o74G8cBwSnoSwJKBissKLny6xnJAqqBxo/NQsFdYzock0MVIpK7LnQ0
xB/oRuwo74ZBUTgop8DDDxLNQNelm9lbNk8hbtXCXZ48gCm+7vR81fCZXaoF8+242MVOhoeWsltJ
XGq2LN+xEig0HWutu7D3hXS4tOlZtO5hlsZlJQK2u0XgN/k5XNNC55wvu6pluCaAooj4AKzdCI2U
NLFnGZ2Ts38U2dQ+gFtxjb78B0wD2YVTC7ijWYNEbQwvU/+W2InD3kxL3qdm1NA2CZh5hxOugWjU
MABHYAI908S5XvJEZ8O5BJTUU6aj+GynPvuE5CXAWOCRpLTUEbkJSg6frcw3pyl/QPg2UeWsSryH
1SSi6QBe+zdDbYybl4keMGyexZe6CcPRAk5LL4hrJ2dp9FEtM/ZQvCT2uha6wq7c79y1ZrL1EhRL
N9sUfjCVA0tkYLd8n4HShlhYrESC50698CETWHONb803qHwr23rab0L+Qt7O7WwRVXHZMuY+/h9m
y73ZKkogRjX1QsFbiX3Br0Bh+tiAK8tXhwQMZIk4Zfab0gpBZmlIt8bho/EbOBNZgzS8x4GFLjEF
bnDpZFBPzfTQIN0I85dj+o4zbhna4qWyDUtyu8Dp4iMBlvWEG2TQJoG/XjZDq8DNSFLXSL0oSIyP
lsU3nye1zC69qerq0ZtQYcrUugazlHka8/jFqx3c01Mw6FImEnWnyRjVI3Rqo06rEKXYS2MYrCr7
QImuctgfSYM/sdyU/WOtZpLg2MPeo+L4UsaK8k664Qml5ux+Khz+p695ujaE3MqrTRKlrGJJzTSc
fFp06g0zWyCqmWcP+E2v/CY17iUB9RoDE2qtZOTuVxCaGCTFFu5O2yLZ5d+QuAzNFvYVc9fE/EDJ
QhxsyB/5ZrrYNBx8voydVhpSk5UOOAJoo9CPxfXbR+nv/ZD7dK9bo6XOesClO+lgPFRJ1BZrcM6i
v7R0gPhnP11cqFB6dn21Y7AcYk4gECuM0V/kjXk5O0E7HMyPVAAL5qWgjB0Zv30vVwcxsY1AAhN7
oZZOesg+Q75wAoP8PGiFH+ptVrJCuVCFb4uQJWFZBAl+lFRVU4AQJH38Ac1IhIylJvcfD+7wCtaw
BJRjO+Q9J3xqbB2su9i5K2ig25Z+ge0wq3n5BYLrP42b1o7Ie8IU/wUyMdh1DupFxTDCvJ9pLc4B
76fiVMfWPbKe4rQccxjmtafibvQnxsOphZ36IMnKCj/JkvX7pTMmhGgT1OfbtK6wYMuyQnIY4vOG
N4k8bIakflZ5I0/YtKPwPWAJm36HdaZUD6dV7YcJJNL7gZcniI8Jzvi+75b4Cxguot+Rd8KSej9b
i+gqiDzlC9fGXA+h4icnEFxi0PGoVrEnOCU+RrWZBDl6YFZ5bUAJymHh6BOto0nRFZL9qNqlSstP
+T8P6qbrR020hA9ITGqD0tkUNMCxn3ngDYWnc0aAfyxVrhh6bYuNbVlCC4CupxnPubikmOOW+0IE
34fJxpkkEJnivUzwL0n8siy7g5H6wQ7aRvbv+7lJeot/rcfTooL7fyn4ObqnZLKa4Q0fK7H206G/
F4nIkpsEPCnF9JN5Prh+I7At/cfYJFOZp0b8z5sE7rbMWqGD2S6caKRiT3qXZrtn2QByvscotQN3
XGsZgDeT2VA68O7hPBBzMCzn71l5z8nl2Fc6ZL2YC5NLubfGIZuIXxRCKMpit68jRQKFlIvnjC2C
F7wKr1bpobE1lLFeCMYSuVD2pSUtHzkn3h9mFCSyhUubzlrlKm92uY/yz2X9sZ+NErIbZsPX5aVm
nDL9uYJl+DaRqYhOc791JjIQ22geYmcc1mP9TIlCmAjVgZ+sBSvhr4DmhWYpM10I3G1m67LhVn27
0owxMqxTxiV8JALqDs+2DzHipfzKcLOmJLlkmqXC0BdUA6+aKgZNpPeH3dPD7h/M0Zlxwh/oIZ0U
qlccwiefBqGM36KPVNpXrOz3N7hyOWeqEf6iHLS1VS++6mK3UWyPSHKn0eNvNpn+xhgqZGe4Oz2A
5wlUBFPA36JL/KlwkEHxtyULnQ7I4/T9EHNQKARzOk2wLnYQf5E1+BmLsWek1bWXaB1LL6vptTPP
UumETtOtjLNB+Rjzr30y2KxjCcKLVAXhZ4WgunDNScMeZqoiXbObbCxcm2QWPP4VgiHrKDfvZJdo
DcLXq+S74laudEn729o+BegLQLFi2hNqeVQxANszi6LS8VhfFHKenVFaSs+xeLmXSIpY4wL+LlPO
dxbnnAhZfIbmE/PVRa7L6L/LeEC+J8H+BpblDGpeF0Fa/4cQferfHnEWxbaF1ifgeu0DtmQg9yph
039BzzNQnEZv6xQ9kMnzaKlU8AieBHnAv4m0vPehucTUFbQKhE1HwKueuq9bfqGR6tOSMShTLd0R
+tSXAiR3fXIM0YDPm9Mk0RiXAi+UhMweaFu2cdtKB5jvIFMf+g3GOcgZkulO2gsoitfJX4/DXLPp
a7bQZaBozfszUtVh1owThLDNwNj1h3bQXT2fuQqADIlDZ/2dI8SSfOZoeTaz9dsyz9tWD2dl8sJi
adIsIEEQuInxd6yAsht/onE3a18N1Moz5m19KEtUX4JNyq64XKe4fcq1Lf8F0HwEMgkTsuQR0R5F
Fnc7C2gYcEFr+Er+NkqPEI/ebhGh2amu5eDn/r9Dvmn+RZroJD0yMoihuHhRRbbXg5T6uI4Vp+uU
GqB1NUVTV/VDCNDgHHBftMxpTqDTM94maG/kzwtYWLb0mMiRSDXHxsE+1lMwsJZEnlqYCiEEx6DM
ou6KMLrrwjmsC5p+YgMrkg/TNIV7xPLfIkQuoUuuyfL05fnjl/7sQTrD8ERzOO6SpVZpGU1vgUer
PmBa8OxHeuvYSew/YHupAaphRAiaxJcDsd+whQOD8tZjaQnAIsUUDAYPCd0U0lF5xJaULdOmWnvd
umtbDfoJRjs6sWvaS8GgoIY9Tnx4+AXlxsJOQr4zv1/Skj5ezFdO/sAdGXNFcnAvA1evkVfKe1dX
IlXgNBI48N4n9D0pVj/yo9fmwE6s/6gR1m2Qftlu5+JbVUBeNy2e0sOZnnQcIU0FPoPYZTKt7Ytp
CugiubSs118cbGOdeNTHIEUjCxp8amBNvjDISZpZ1IRPzXrslfaTeoGKIWHoNL3fRjSYQZr4lufY
VNHyE/1VRAmAHFPgbL0lRuUPPaRfulJM4KVlxZWTrpQKcsNKhmLpEMcqcD4acYLWOnpbqLstfj7A
NZMk0NjJuvE1r05FyulUCa6Y7fDL/vkJbJOJWC48SI82qu9mZiRUy3K3K/n2YZzwcXU3f049ebPN
Ixz4XsYHqPJITxvHpmOePuq2pNNxQBrvH9+UB/bencGX+sOA54xhJd23uVxUttlra2o2GW/yklFN
Z3LLJ13q3gGlF6Z8f203FsPnp3CILzR6Et7FnDW+8+91On7J8LFiDnVHE4PlZ+i2QNpu1NPgw/70
XrmxNsNzkaoxMhuEqVmYErtQ9AGkv2aq+z0sqMzzhjASmTiWnuGkCfSasDgsA/PPd6V3xKU2s7AD
6Gae2eEtoV6hi1s0ogqAQq/+2IbhjlOruvmgn26BfXZEyJB3e2v13bJ0aR5UyeaBj6gpMc97BkEx
eobQ2F3M6I67WK/DfXmpl2W+OiXckBuxgD8ZUDQNJ/TWTgGtdiNnYlFZqprOt0OOw18hG6Pyz161
V2K7IVX2qI1gczkh35vMUsqXv3JIrZ3RaAfBfbtewsUVArxcjpEwhFgvmyP1G61IPPhF72PqN9W3
WRmBjVxscrHA9U2+rSnErbNjJrz/wPcIiEPmTQs9oU2/EikHBbM5SnDiWbsGi/XKl++HjXEblMSJ
5jpmvXaoGtBQ47i6RHN2QrbZAFpoBi4lMJn3CoTHXpAEFv2rGK5edhBx2n/dHORhoCJiv23HFc5o
WZFy/oPxJFUc8YXvjn/OYTx0f/yIyxzGM9XmF5Lh49c72PbCf9Yl8z1bVXAPS2Y7oYIqmiEVWoVf
8ox6moAGvPAWMD4sMev4lG5mLr5JQKDSuqsRJ92IeMdUdBNstmwXhmkcbP3aNqX/ULJP7aWjtI+Z
ZyGbiJdDHoXuUqDbJ9NCgArliMLhl9jnBXJArQn9L0Z1vAuMRvvVmDEsGBKjMr1SGhdFUbM1Tn6h
8teWStADG15pT05sglII3FTgqQqPp99AtJT91j3qzk66oqzXWmA7rcBJ2+voHLIxLTEZAE8mv0//
y1eYjmnNswgELxaU4WUVlsILjKo5gLtE0J0Mv0DuszdhazdPiE2/0Yv3S5pBZA5oYkt6ykrpyPio
oXDNKOc+Ok1e1jOL46ih56qlM0nilY2yN5cnIaciVd+XoZr24eTM0SFUbLr6qs2q4bohlU/wdPkE
TAkkAaCd3l05bup1MlXQ1R+c/geBXZ/x5v2U0sMtIxCQJ/rTgimoAlsYF6l4cuS5F8L1HKDR/1ML
2xFNOzYFO4Pi/l64lS+YVBB1RUy+fUsxIgDfs5dzwmJNBR63gH2jQXkT4sVTWHNPXKS1FcMTHZCX
jMnmf7lVLZzzS5cQCCWck2zmNGnbQu+SFGsM/rURbA8Q1V33NOrhIQ/5gbkl2PegBiZl0zUs1xan
z9wewlul/zryU4ZKo2yAqGrHASDLB7g7dyfiZBB+9nvkZ0Pf4/WRoLvSmuSybldMfqYOnCXHAAsB
wVbTo57UbFOGGSPm9/Tl7uKYLkh3qQ/c7Rg3shD50Puow7mO/iZOrmFxZ69m9OrIB6YYp/F+jNha
9TQ8oCu9RAgrhVcJMRKpkFRhgnrJUYHyZlU3PO+3vf1F77FKrjFF7J9g+3a3heuBdxMHkjNXQ3P4
gO9IamrgmSGkuIBJv+xCj38bM7qq90PIL7EgSXiq+MkMRDhGFIFsBrkYjogsOtqgKMVMNr5vwtSX
TAkKFvFyNKzJvBitqxsXX1yxhB7WzgdqhwlwngeXVYWyFBrky2q2c8iUdwBLEntN6Lt9kt/hfhLE
MWFH5hhHPoC9bMg/kvNiOcfxAY10eNwZpFDnnKovuT90mGsPOh4JmtQAKEsC540kdwJUIasbPUcM
Z2d/rf6agkyIJZp23YED8kWLxGaKI2Cz1HCXfWKCjfKTHeNQOE6rAVfOUEl2703dk9Lr+Lim7dl0
UTTtRyc8z3n5nBvMEL1QTFxrgogFwmq1v5NXDXgtPRwwCGgUJujCJFjASYyw8po3DYPr4g273xR6
hZGMJnFVl4TKlx5oKFVg+x8xpW1xzPRgBIEgUH28ZBdCXYv0LhR6jKEs1w1zp5QU0VxRlSsvaqnP
ac+aXbBlOjMDqz28cOU+5Tx1s5qTQq87pEIgXRAO1i7sV5BwsvtdXwdwD0FGcAAM/1uPh/gfkazf
AMyojXPmpD8qISag0H8ztnkx7khzJObAa67SqVr4hnVCQakbkMRKxmirtr3HG/2h/70u/p6kqB2C
cGOzPyApn3SXyZIHF+oidTeSEhy4aYFWXJDnvnKHtpEzOG+YkrsrP+3n/w5birBeIvoA/2c6a/lg
wILlNg3AR0GtE1fhrDjyDv90sHPLU8vbhz1FIIBuUQl/W47JmOzvB4rl0YTBXv7H9+2pryJHaQHU
W9lJhCgNcSCxDOzQY0O5kBWztaMArUcY/52c1fxEHWJqxYDyLOJ9sAg5Qw2FK0xEy9fpU//hG2gK
F21BZKOFUISrt2hqlVQd1yeFyc2lq1ndHRvEwoMFXKJJjv6TnFvn18vA/aFXM4uKRPaIgco934YW
NGAt7/utIl0J8Tje7lx0Ud0D9GW7YK2FYHGGnGZXJsAHSffFwgE76QwnD8Px89wzCZt8ZNjhuVn2
kJWKMPwt57wHyaYVVH1AJMyAJM5Im8ukjiWa/jfvyx8YtGPEQKO3Z+vRtbQyJu5i/vZ7MAbQrgBj
z/GVUzY6xU0SsjPVUcw82LaCyryRtQoqc6npxlhf6i5gdCS9e9jGa8ELwJb0BB06sYEkJFc7kVx1
01R6XlugLiSlbvgVfZjpRGGKZ1g2ADb1XlXomZZOJi07ERSBwlp1FYHrIAkYb7wAk6FFzh/qJquL
z9jV+nqhhY4uZPGc7zr7S15I/56BB1RuLvyxP7wzWD569ek+jEvQNCJjsVHlmJrAe1i4bzi3kytz
71nhT0AYUrVGwXMyEQteg9nHyXithG6IF3OCTIWH/xJwSFX4kyoWdHfI/n6Cwr3Zf3HHm1TsKuKq
K8pWa3mbaHe8TojGVQoICBXqNhPWXusxjanaUADJ9Wsi4REMgpidfP/YNJ6Cygs3GmsiZEq4vh+k
QZYeSq+e6p0OLWH39lcrSY6r7berCflY1xnFdgBL/YiNQbUtLvmhNA+mTSOLLiCfE8JxWpK3t3qg
p7rt0kvEpEioPaxvJbi5/QzDOvYDdBWMVBmELwsYUqJnsq2vRt7GT6cTcEVRQQDtJQHMAzjiiXaH
DUca1Kn8mmOW+Dc/s0a/Eq5xHGR0P2I4kQM9J+mLcyXp7/7T7MxqzcQACHM+kg6ZWEQPuuJ8AiS8
rN5ikG3VAICiil0aJBi5fKnTDOL80q3NaMwYB7frNy8M9bYDWq+7FH+smnW7SDlLrX9iKN9AU2C1
lgzY7F0MBwUTBuUxe/q95BtLxpGBdtFr/y2OZeUWaufB6ATLUdJoyLOafhdUAZGxVGA1p/RZZv9f
TNWMuKc/O3Cv8ZXWiuOYINU5l7z/zc8ze7Nu8BtVdt37WlOEqXd/FU/6tOHDcjDfL4Bp+GKxPgpY
Hi/Fk7cINj2FmKLI9CFRRq9GHOSv4UBlSk/7QtrhelExhaQ0qMOKzM9I2Aenth6R0d5JpQIBzjTG
WMqskSqSvqsmoi1GoOUJ6l72QmdUn+QnFSxHiXCHIojDGfhBWPIA+LpIStk2Oh4XnFOmW6yFGlnk
QKE637QO4mcSJFRyKiUW4+mDgO4GlpDpWZA026a03X3F+bHK8WekyHixoj+3XZehdtKv7yTQRsL2
HpEE8MkKMXogOFBJ4gzUQb9JV1C2XoNMP25aZTzqK64MloKMtrWlAdA+0Pmh4cBhS5gueYdEXgtk
8kp9Sed3Av+iTZfOfSe02uSCgyNlOxqBj0GCzJkoG7FoDAzYOE0MCsIiUYfgscDHzY2uzSHKWmml
re678cMZB3LMiEH/zJaq/rxmFEiSlAbp6ckHXjcstwouPJXMpMm+zZDt5WsDPRAg2IQsygJrqayE
6EPIl/5T1CyFywJ8F04MvYsSvZ/eLH/nvbSlX5wE0nNnF3yFzOOTpJ86IchaLQaqYLhymQB6RGre
gR6sgHlOHlJM0d6FEu2b3qV9nOmHxLal+EwTQWsgKDUa2uy+5bC/5OGSd0/dVNgFxx8eM2Wv78TP
lZaCy/nmp32rGUBn6JE6qI3CaWlT9MqZXc2JvS4s7NKhbZrwVA0cEumY+lG6BbUhmAet/PCA8DJi
gXNDzf4QWoQ/437Ei+gyDBcmSRuzzFTMzNxkNFFnFMf6bpVASCDAKeJrhLaMXY9507+9GwzJdKb/
sb9kPhO97T8EtrbPbZIiRl/Uso8Zq3490kgdefe2Ejb4cACD+2wqoDROVgorlwbsDj1olYG7qeeF
hVNEZQi0f5hWh4pHCzeGXl14VkvYfEI7V+jMU/xfBbI6xjVKemnRBZKkd+pUt+M46ZLvJHT/IuGD
WXVhQEGVuKb6+9DeXOs5BUmpVefcShuw5l1pUCR94nW+WPAJRiz9+aoIMNtTY+Akel0yYEvlwC3q
UQPQChERo7qjrIe9RrUkQ00QS3MBwWNLnnD1ZTREahAJVH8GVVriNy0xi9Vu0pwV2ITr8dD3WZUQ
r0Ly/qUAq4UJSGrE0hSduWP8LjP7C/U5iyWt7SJzTT0G04h2E7zpppOkQHMDz542onPbjwjGTca8
j9tfps/X7JHPzhzPcwP3upu6meTmR61cqAdDSsCBU1DskNCVbumE28jM4L/pDNZiwq3rBsXw1JUr
DbvEG5mmnMaojcrAykcc3zLmmeIBzjwHjLqbh8eQEZfoQd92k9gP7lqY2GgZJ2lCfJPhqV3nAS8j
kAN+4ax5Sv0NN8WxYcCQRcFObQmn66JRhtkqOzeS2dpFVrYGkDR2UKX9zQJdy20Lb5qKUeimuOct
WrhMNu14TNRa8EsO8xCQH1DGEd8RCRpSytaLrBmI+JmYea0L3Ddar3+hkXC5ZgIMS66pElKIjEzb
ZhG5UqI2XCITqaNS5W5vE/EmirJ3gThi+DTcSbKVuZvD0zaa5lSwG6JJIksG896g7LJOhxb0N53+
7Vn7rTXVatxkCUQVkjmevxqOo1c+u4C/fNZl1C+YqSllM3mn+OWjJ8t4mtiQSi5jX3GU681NkInR
NfGGbQ4KxwUFMeQhdng3xEooG3g4f//RGKerblTaRJ3cUK0Ci8+NV1M4ePbKaoGl4qHpHTYpiR18
0X/hRVubdMq9OMhWeD6JyL+z8cGMfNaiV1GMkXlFDp+LpGQyOptRd/EbNiYyBtRfn2yXAMrH7Z6D
W48HCkUsUibVsIKFLTzCYHPqsE35Zs7g5KfefirHnvgSJ9nhu5iDEFttIyL7WAsIEfYJqWE3Hney
5OrMrC8XUgyRt0+LGsT3bZHqFaKPxSsI77b1HtClVdMRZ0coOnQgGY3fyg4tlcGq7UI2IwVJ7YoX
i7JdA6p8S8lBOEx5MUplVJDFZrUwRYneZEyn8z5gOMiWFd7hugMtUYZ0PrMcRTAJqCXSLySwrxpr
2u9/1LwXXrH0T+wzenh4oazLMTWfDk9yhUcqIKOisMf9aovlGbubyZ5U/nEOdCEMzTH8HAWxxd58
OQBMOcjg+eGi0Nm8aghrGivE1jCrPUHQNEmgkHTq03suzyhU8KxpWLtzVE5oDNes23F9HTrkYk61
Csh3mjN7ESeBt3zBygGhpU45FsLHg++ofY5Q8E1siarlMHE5xpQL69Mt1/i0opUth5NLPkSf/o9I
adsEpVBr29c1G5fYCrOpJjMGFfRADVx9DjOE4IfizmgJArGy81jQVgPLnEGjmqvqRsly9JpjkV3N
7sdMFuctIbU5iLiRySXHOTdK8kzMNDUvBZFJfl7fGuDmo1XUgG06lZfI/nSERmM7Pp3LJ4lQ9K65
ZntpXDQZAGMQCftLlosORl6OZY88AABBSbzm7LNFjvBBq0TX2Mux5SV5Zt639ifWypzo270NlWkI
/oqL3JruirZEeFvdre2bSNCRJwDOWOmWZ75OVfUtmW1RxNFJmfdhrn3n97Gxkh9wYA2ecQvxmY6a
X4ZybUDRg9swqKaSZmas53OlwiNx+wrjZaI7US4QNfIrm3snYl1xFbPHf+vyecv+tQnZMYxdh4Gq
/HwptBqSRnFBUcS1qWTlI/dSGW/RilPXIMot7U+/VWjmMfYNqcxQPn6Y+YYUL7qh43Ge3SRAsRj/
bLgI+JC73j/izVZPFSEBs3NjsDKqb84DSFmRg52MqAJR3yIlbKfRwzzGRHs1IcNuRZ5/nZyPut2Z
0Z5QXKisOKCC7p3DoONf2lQLRWxxWQgGF45+KIC8liEDJYIKdMy8gC1R0qw13RwKyoNFt5dNxMt2
56QXqkUvaVNzwCeagpw+giDctUcGALPGE4x7wXD7ogQxgLzRctJrzCOJGrDXP4WPxoHJI0YEAps7
IlQZCu1K//Y/q3BWaD/nHYBG7dieIwpO2akooyhukjWG1gqdImrHNRzT+nlHg8IzEa2jtYijBZaA
Ix6sF1B4AMq99IaK6nndWygrByLifwzKafgS+JM3HR51Xdwe3p933s8LJ6JyRUkj4qHipXw/05MQ
pPXwq4+ticWAbWt4Fpc7INqMRwMlhQX0YkPtBKox15RNykohOuiJdJIwQ87f2HSXUhO8UMIQMoQG
HJlyrYZrUJHuhN4blJWQMAvfb8bA7naQCyCUwIWnq0FHAGy0PuMV0OqhBgEdQgLG62djjdzgNu75
EGna/N4exyUYKMR4JSDATl95KAVXwjAqucwBFVmgruYZTQwtxHxN6Qxy6hBsw4dSrCfm1JLBz7wl
gV5efcff+1HAenJmEg22x7tlrn7cNeU0JK3laLYQE2riSITJcPWqpJGs35euoXBjoyeMHv2ytraR
hEzZGFq9nHce6oV6V1ngAeZjO1eFGvUTJkyWcECAMOKdl8J6RUM5ixC5HggeTCywCKXyPveylGFd
834/ZFCi8Roy+zMHK9Ps2hcGWURy3BbayO0GyrAGno0gXvO6vaxRIzn2n9uD0aWBBCHliozFjB2n
YVWs8mT8qdjS9xEJ5EkU4LMb7qgSC53zhZcKjuc+LNlYDtsdOaUO3/5Lx6F5IASvDJWZiNS33OIH
9tTs+9ZKAo1kqcyayNdeMb3+OHRd+jq+g6xstWFGAbmhGZylJ3Cn7XbpQux4IhdUF60NK4WHhcED
eCaWFqhAA5CEx6hBdceU4kwrT97nqk2wGRHhabmzZ8TfBukk9JuhkOg81GMlwgNcdqczkedEYlZ6
s18JVFIsGO+ahmqh0w4fD5sjMQ1UIaZBLm7A95/G4Lsa96o0MYWV1OZ1iFRMGlycnMh0J30j7q7d
NTmVec+yw9l7sALKqIqYF+jLZgZZ8D+ZJ6gcjzpUOZ6OPk167rUS4kitZk0iE4M5Ne3wSBx3SmRF
gnyQ8cnMFNIpWTLKj31p936RpzOli5kqWB5RVynKb1qK1bEAgefYlJSxUKS1qArSg0bS3am4k6bY
p11e47LHZmJ+aXBLfubQlzGrIIKHyG2Rpqi57f4iWHalcLYp1REuFdB1WYQ0Cuw12u1GNQz4V9MS
WPns3Or3a8OuQdC2Ej2p/cgBNf/Z4giwvT6kxiAwwxCYhMBnxFVuvKDVX40rn3WQ/GgVAgGRRYgP
KgvX8X+1MXQ4KWpKDIvrJT6QZrPcP9nEucKCbyMJP6UxFUmGtserDwqY0VsbgVRA5WtLMSMH4gNo
RHwhgntnbIGKujGcp4EWmJY3UE4TNArcda+u+LsJ5cDu1v1lh2hzWZhK8Fs82Phv7P9LTCEPCi+H
/LdA8S8p5/tBZaRMnnI+elBisb0viiVm1eLishW6au/AJIscW0hp/Z78dyVGnW1czux8gb5PBmUr
G7MIZ1919B59c9ithdSUOoSBTSrM1waRgLfa2hCxF4qe4ibKk9wzwgBsvZDb9/cXfgkeh+hbEJQC
U7fWZzonhehHEPKYRXPeTLirmZhY464KU0tVXCJIAc/cUM5p7I1+HzIkOLwutEYRnbEePnHV5WkC
T4MIoZKpaAvcCjuC+PdkX07Vf+oLCxc6MgLYxkGCvA510v05xRSmD7jq5kGIJlrAnIhybtf7VrGr
dGi9zE4lZTjXQ14qYBBfoTJo7yFpoFCM+WaIhCZkcBfhMGc6fx15lgVP/ZCKB6TZsvU0LZmqAJ+R
Ue+aP48L2NStYrofdSeiEzl3nXPlHEDEa2HDY6nzkI6BSCFyKmSFpghf7sUEyAjkcFLVfu1/xOUX
ZTMUVq6jWnb4TwBVIOpLfLaFciVUeVzQ0m47D7Kfz1Gw8sP836EqMHI09zTrh7Hf4VW1aZIFMg/C
sss+WPp3Jble8PK7e4BeUsr2mRscyVu+RYbgP3uZeYMnKSWV/QwQHsTbhZrNLbJrkQ7IZ4fh68ir
s86DjiKSg1ovWjjYlNg4TJKSa+qcvqdO9Vea7w0E5vvJepRGANzDmeLnAGwi54brKRPsiPILhJDg
GDkq+FsAHOE/yvWXHcE+KZoRvZO4YRUqe8aKm5VJfmeamTfvIA9F/sJqGtoD+eYkuDWuYJEjk+nM
B6UReS1MLO+X4/jTKabNghCuc+gusVvTgmt3LrNJb5VEqkqGXDMb7wDuvvGvUhrIn7IGcq6r4lCi
kDnHxnwxIKZXjR57MBF+tNMPHx2SOvPgtBAk/Te9oE1cNQYwpWb5kz+op79Jf4YumWQ9nKcoGA17
N3Kzq1Ym2fS6u7WLYpJ5tdDGdQHIAtlURfPOPQ0DrTPziCwK7YzBf5vjM9HSAQleLzTOTcGVA8Tp
xjdPqTqk+rjSVr0XdxFWx8XwGMQfFEqOAjqshoGnDLU2wsOIwebImu05tmlNn9C1xWGr4cBZnt7Z
F9aZh08Pw3SNi5HxMUp6h6Btp9Y0vtwm3xD6O6q5HjzK+Cm/BlSZxYd6+XVpnk16THlIOskCYGIa
zyg3ybccFKB5PWMawnaJFHvLzew5onnSRfH25sbj/eZMtmKmVZFQymbZRIFC7zVuuNJFIhwA6IBI
6YKthcy87oY0S1JSARmMPqXM3y6BXoApjQbON5MlvMIGxH5CtpyTOfo5LsPm4zOWpm1yCQCbLnPR
Vgjx3E5Bt9tbf8CJI8Igdql1xczDnBYvj4EaeGWrU6ymuwcuPmbPEnWTB4stxBlTvceViw6J5bfq
RLLAMRuyItrscofgRSCf6sdq5g/fTZyOGXt1AhMPRcMjplWiu+GoW9o88kLJgN8tq+FOR9yGN4eK
vnMbfhc27UpVD/+1TtdIIjXv7CBRwM9ixT+PV+DgRe9fzBuK3tP6Xc8uYtDSfeBw68tyo8m5b9QL
CNCNLXKc1nUw4lnQWzlnVWcWzoR+GygZDtm/RbgFcVJAfeX+lKq5zp5W7mxKAIN4klNxxkGxqOD4
asFZ/PITq4qMDQIbCAbKFoks33OklLS/eMbWp1GtbHYJ8hkAuOKTqbi8yobkpCi1Z+jfDQZB8PQg
/BpNM3bjdsTOg3Nw21ZcD2G+izz0k1NdAfQVTm8muFZLel/BdpLTCML+yHoqrxUyPL5ymRGwCOkI
ubrT4W+HGI1ZCP3XRugUgbYb7N1gTUFoFM/1YFvB0jGZNXMicBsGSW/t03hqyAYqlv2PwpsWveHg
VFeuu6zkqZ4DMPNiVfD97HH4lotw7ayFKqfPtUgs3um9/y7GNHvm1Jx+39LpYXHpFUMjSKL5j8Sa
EGgz43sswx94Q/+waTom2fkBclJq4WsakHtSF/COx+21nzAhBJ2Bas8xvEbtBA2hoNVRe/AMMaBF
k3ZsebA+Aibgx/Aj68MAtPrzcs4quDh/OTM+dOz7cD/R5O4WOU+dFUuwZzDD7/diRVjeTjugKAf+
tX/g6nSVe9cvKaUNXv0/MHE7EkDbAIyu/OYdJiTg2rXH5qoGuYbyqDjkUkqKP6InQlwqFEqg3tQO
jnsfDV1aNIWS75NfKcm/g0raPaL+YhaMuk2ZvkSrt0tCBh6Oa1xOr4+2hF2zZZnlc8fkLnv42A0A
HlA1zBYDThTtCnSZUY9fZg0yKn1KW4DJNshM23j6DYFQW30c0Fh2FFOT6JWY80A/dNRqn5T1Lmal
y0skIWeKrtN2lZxK+qp6rdey+44pz/+m5qiazx5lZqpxVB20efOtLkmyUKOicjGEl8wyD5gD4a5u
vznzizIZRgZxbWoeAuyY0wdqyK+Wq5+d6doETvzEYc6TZ7qBd7ZC24OU+D0XSIh+X8isq2AO6aVA
soLyxJyapjeoDlwGFxoWkjiPSw5Hfz0O+r734pNMvfzpPobzeAdC0ptUdVUPXA2iuZy5erkisBTC
0FQzUr8nCcm7bSYRoIcqKrokvcA7V9/7Nd21wxiacDBMWqxgdT5jJMGtnwyLeawsgL3S/7pqKTz7
XPWQ4h8aYZ7yMIQobPksodiO/b+PmV+lWOeRyM6lxgrFrly1s0TtyWcOtIbSwRPvWRuzjij0ppPH
GwVRWhD0EnGHA4/kLBohBK/EYQCw0ZkFTxsr0PpDxPAPe9+Mdk+3u2mp8L3vBSoJob5UromF3Qnj
nKwOJ5PVJXvgSCeSOS+ciUDJmcILbGdrjrWuUGyXA8ypaq/r7TOWFHOZeAEbPP3UszngbNEj73gF
qB0mk/rgH2RIen5sf96vXp0w8FFMEuT7C7bbmNnQYjBqyycMdyQerL4EHEgAnJZ30vACc7va/UuW
OajQ5OAZ5mPzQUXhxPkkew4XF4nbiwwTcgGETlZX6uqj3QRUvxqfV+jmTtiTxnHQTUnEAA1Uc9n8
1YtaWk0ZHiE4/DLZ8PlvRo8Wumc3yuamIigCOroT+1VoO/cvxVLWT17zNkVTF8fcUJUSJEU0HSfg
f/bJQlcFFlBq5Wr5NMMy7A3wFoFqVzaOMh88jp2rih91j5KNUXBAd1PvnpW9ZQn45VlIeQISHmuW
h2t2zyVz8J5/juRKiBc7An62p7TgL6xsY3UEQut7JHoFRaOUyak2+rKQstdoAz200nkSbK8gnkKk
+UOdVC5T1Pmyg991ORSJE4fIISEAzzVDj1aY83436054yxhkMC5O4nipTbrEEKFq2WBZNa41WcQm
fD95hI8cyZNw5jph23DET79kttfLyJrpQrBRlddjWxblIgVa4nhanhqCV+20+zg8003U78lA0x/Q
ivJGHS+9awBOQ/mDoq1K5X8iMq9U/Wc0/sTGGP9XAS32bw8Iz3oH+8rSoI7YLhuaRLChduD15fLp
+lsAvnJ19eTjC1iGV3yuNEokUsctQif1ZkqQxPatHnKUQa8QpE0/S0zitxvlG8eRQhCg2T0Rzbay
6zk2HrPz70dtQtlzNh7l07cYWn1JmQb9BnOW6fyHfxFGflMe1E1nYtsMlEuPb+X2kVij3cq/DVXI
Enh6Pvxv9XYrWSFowJcG74D0BbeZdWciqg4J9FMozmvZpXJvYo1trBuCSAvh36TNPplbK6mLcq5o
sRU8fNcuLX0pKhlp2m+1Ly5DRdQBL3j6giV1hVW5BNcSXzrMb2DWCkCvcMAgCw0SXKQzWO66ycdG
sZCFRytZJLeqc+XK3Kw3wX3IsvRs85FXRIxd7NKmUKXx6nk/kdzDH60D944mccxqRFu3JF3eenfj
MxeSAmzV2EeY2r+jCM0mWCrsrnugaGlzwJ/iW2sHR1j4sQl55ZvhhsPqa+dgCeH/TwvSTy6/fFH9
mbzmXfVSPeKossskK6Z1Ayo9tgpE+p2tBiAQRjkuJdyK1BI0OBkj/KivoxrYWQ3FjtPiTrgbBZQM
rUsKhekiFinX2LbEJAWkishV3NxOgy14VSoUcwZzz6hW0no9NUt/PBCbaz9NUdSCyJIzxIS9u50K
2r1wF+6aEk70/DZN40QNPgEr8mI/9gn8H/ZEN8qJM90I9sZXxLyGjCvojS8lJxcyGIgszO+fjwRQ
e+jNSYi4LmYQ14n+JXXWyCgx2ytDDtPfOT5h8VC25rUWZhvoGDkaRLt8eoIhxpMrbhvgOHIi1a7p
3HSp+BGeVyxg2U4hiZJP5ZMJrRb//eXZ02Sepv2Ben5QKHtHY0NK7jnewnOcFi16bPZTpyInCj2+
QZAGu/AgqiZglqT9Urs53C6MVYlkr8qGupK34otD5w6p9KRX3O1k0GSIsvHdWIhS37wmsS//I8WH
2VBuH5mKG4Ksb6qebvBZwG5PsKKATQORY+5NhbKzZFiE4VdYTssymawsB6mK7IUdWLWM+fyBMXuw
2/T2wSATOgLJjP7bBses6GYzgQBlGjNDQGIIljr8YcZLsDc5x3ondYr9XH8akmHqTky7JqPUo/Kr
+qKeusdvmdq48i4wFs5dd3uaUPz+yshSggBWfjCVSZxxWreTP4TmAIUoNFTyzaamL2YBA7gqeR+X
8XWKHpLj7syUwAo7wt4u6SoNcm6FBs18DZYOONFORTRiaWhydRWi6z1Lbl5XpD20hs6JUu+g/DEm
WW/3Bt0suBcIqXWcsg0saZyiJtIllLesB1BwRepHJPyBcfnrCt8oxPNlln/TxX8Wx6MDjaE2UwZ4
qLWM/xdwEoAltpHbwtPQ4UWH5p932rJLZqkXFByDoLEUGMI8tar9EWLwgJw82BahKTM/XEyAbTTb
cM8colJY4NslhJDm18vkGybw9cPR3AughkbEFzuwckCyRC2xel6nSJk1CnzQ7w+3V6FssOup478Q
0B/0EgEq+RlVlDHoLnwOJwsBMG0Iub8iSmPz2rX+qbzcotBoKyXaqyNlCcVBzPKBmd261nlscoI4
2QMhd9wrqIogtyx322Pf0be4zupGVqm4VjC+yTCCikTyxXgkLF8bajcD5/Fy1c/GBpNSvezaX7dF
07KimdHyX9KSsLPAGNCR1JRybU10PTU6ULnJeAjFHX/ud68C41qfflprTW1foTdear+bwjjiOwWa
gb1/sVl+fm34azvTTgk3yVyg5Ym7JHe71gRfikRu5X/sry2s0flZHF495I58eyKyzfz7xoDNN1xu
wnrbeNiSwqG2aHDv8++bIGOHiVCR9Lq2O59It7y5UIBBC4dpY6Dy8S3bjH1W5+KYcuI15jj6JoEF
BKFUP45NKcJL19KzAlVpcoc9oxNlx1p7nm1nCz8NPxV3NEVHSCRcJWmpUx374YUstpGlp+A9BZZC
kwNz9MKOVfy0OFhxTa4tyCA8+XKYTkjsOUV9U1qDokSCPyPKEJzYejgxrgQJoeByPr0BIIoV6V/9
i50UZP/NqCjldemzTLqwG1KEFSFpuT2xWR9HOe9rJzC6HZZd20BPJr09FbTU+x00ItWwFHHI0ufE
vPARGwyyuqjF5dXguECA2+gXUtflbGwHoFvWwQh7aOIz91r0XhLhK5edwc1FfEA8zc4fhEWfgm0T
k9m1eLXEwKHptk5EGYaXJaZ07ilvAGtrxZiPGN1qQP8zp+7znneOGG6D0G6SvVR8WIsVK6iQcWgk
oG2D78qlaNj/ShyV9iCYxue33iRDVaX74drve8gyfU39dwWKk6d6itTw5Xdom8a1LHRuonbvj3CK
B1FonG1Gw2h/iL4iqWmUJmra4NQwy6A5fZn3i+K7JzItQURwHneaKbgBjvbIrYTvLBhFMXFsG27w
xVQInCuvWyC10xCNmvLEIPiOvuA8zmLSJwHhdwDTruDIHonazSgDwFvAQNOnZ3stgDO4uYj6UJbI
/Xe6daRdaEnz+Tu4zIxa8DCHGH+5O3Dq/75Z0f25ml3rSHTUkcpH7SWr4144UBR4vaUdMIP4apLr
ETlwj4Tzh7CGNk6PA92xWFY4+BkYIH9v11+VrQbUjGUaLOVNy83bo4n2JHztVkvQ8CQfx1jZ5Fhu
32jFxS1e6bGmad7rbyVlYoefFN8VPX1RBNNhpVf9uRdkRa9At/KKxWSe6A0iUTRuJT8CWNxVxgEs
WjBuNXWrg0/jKSuTVxgH0Ly1eo7KExO6TCIf+SU4KQfEJZTUAAZtwUWOtdO0qVNs/V2mm5BwNIuv
xhXzWrqfB1TBMgYLsf2fQLTnoLNO843MkXMs13LVd8YeXcK2f5vxKdYWglzggekuT1oliw8W/iG4
h9MS3W52i8vMb3h02ZY2WJp9AAVixyyYJk8VtsvKu2l3g5fzDtG/c2fnchVqF24Goff4bL8aamLX
+rStJ19CZH3C6n1HWbHDLQ8wsBHXseqHWLZ5h4k89EbvYB/uQh3a8mxncGDJe/G+a2LFfbDiHwHV
by1mSYtM9GgthOp8+xZwvkw7/pxyLCr0OYWS8mzo/OsVsCfbp6Zax+STXLKdSyE5CumozAJxb8v8
53XtJpijNki7GDAzQsAcwJTnJ4gJe0ZexrhCu71llbIVKKx5NT19985Gkn3Sc7HOkEhXUdWkALLj
mRPAo0u9i6vf8rzc8q3JKaAVWPv19Nf6uwFffFBkyWKC190j8FnpphkeI7lcz28J/03z8YCr5oJe
jRtAA9zO03Ks41ElBqz9CsOU2LEClWvu6j55jhJk7ud0k8Tv7cC+HH0+AledjPwODW6dBz8hWp5e
au4Tm4LQHKoZk/TMjfV/fVGWbnjK8UX0dfTxN6QP+OrhI9lzWcPUhoCM9pZTLraHWxOGULkYezc+
FMBxCXFTjzuH2ZlKce87JqIFGE7f2iHxhIDyKsvDq9vYhJtDQSu57ZX+IHyjMArpgIezbtxLOQYl
73e0+KREg341dVZIEMBIllewkPOyqDNHHjfi1XP8MWNXS6kT+3R4zbcVt1Z37DLVpIRI8DYra6Zz
iG2d0tuYNy2qyvNv58x71USOhOZ58XnjP9EjgIeyuUJHk7LAyw03uWv5HhnyhuX1k1rDi0/r0/fb
cZNQCYdlea5zBDVY+IUx4ZXAhy4fmpdWH6NhtteHyPu3uIEmXhp3DgElT3pqH7efFUcUMM2pjJee
hR0UeIYWfPbSERL4QsbxxbYUOkG9ukcr8Hy5KmSZf5dRYtKfQW411RxaXJt+ogfW1Aqcwzttdrae
LyNc2YLLQlQ/uqZwm21lTtb03C8cPlebPfp657DJCqVeafEYVLXEnB5MVKWfK7F+eF64yJ/67X3u
7LPKs0ZafaEuLknra0021XciYUpthrSnF8ec8TesPkxWlImYLr33h2O6Evi7J/naFK/AkdeDJqi3
M1cjncEKDV5b4CvWtS6XaqK4EkKOFdNk998rP3KxjMLg2xhgXebPb9vVjvn0NneCp0oNS9DHECgi
rLutIeIjWqROj9o4Zaxegr/nRN9+ohZVi7S6/mf4mCAd0wUajJ/1TONqaDfpqTJQIr675xMo4rRI
R+93xycpFA2GXSyoDk8opTPkZuLbU615xKHkbOjYkyXU07QIx0pCnUwbPlifYvyTxcq5g9feGsY0
g5p3oDznYoqBdVOIpe+Ictew2onQAFvFL4uKbAS8brXde51skaKJxDDYzSW0WDWThiISQD0eioTE
YiSuB0B7j2U2eLTbYJ4H8NYDBxFkzNRLebQ0vkEH8Uy1Ym3svEAuayo2xZzvAvDswxVcUKXkGQdL
X7V/dvbhLfkrMi7WLH0LYgpRXodAGUe5bffedzgy/AiKJ8jc+oOVtPiiRvy7QiQLxGMWzedWqaaa
+4uaXzv+mdXLfW0fDBqPsxxcTCjrZmFjNlN+sdVQYWpgqyQ7QB+XGw2Frz2uV5dO8BetStfD9VT0
E2b9l2/IYByjGRPF8/pH3IrlJNDdh3MiRO7BRzmEz4zdrOvFCEoCHD6Na2XXNJ/wssllV/vcOd2K
QKGwVQBdyxNVJ9Km4HFO20P0Pa5mTTe6yUeoDMajJmnDd3SAwGT4ilyHUhUfYOd4frjqcAkG2uDc
7lZepZ4tiQ+9bo3UKGgwJeaVBtzqH/ZZCgdNb7blYlDoCD4K2WtDmlteHj7wJWJZuElJp0sJKJo2
/hP91LTr9/lBHBdAq4fyC5tHsBip7KckmbB+amX6FDc91dMPuofLqLRco1MPWJh/YN+sR66uKzf0
qRLYNZkYBfcDy3pu1/Ve0N7QR8GeMr+U2waA+eflMtGxA6ilH2VeJ8420QWgianjKMHUxYjHHZ2s
eVoTBCTYUDCz72r35liHKwjRmW51/Fe8NSPS9UlmlmB04+6KRBUX9ZiiXpM8JWeW7nOhvM4OmEsL
nfRXVOxlJvEiZmfz+Z3Mkg/X9OJPT9NWdSgkhNEU26WtoBxWIS6oxL2NQ4+n+wbtf5womCenVmhU
JswrvfCoJHzLmaKLxE2D5t+Gt62SVVIEqFEwPZT2eOld/+CPSp5uL5aginIXwc3QMle4t61lakSS
S9jAAsTFUnsujh/t4utcyuZqU3D4Y16LQ5LtPOlTnMnhvyvM6+oN/40lEm86fddVS3dx2PWuOpj3
xITeGjruVqSI+OOHnKXhqs10wDxI5O8q2GifpvqNjyUi6DodtA9EVUZczOj7ar/1ESlmCZFUGpY/
eor13Cj1Cpt9VTJRh1JUxX0/8qcWX9NCNRbTeoxosk3r6OXVCC6rliojtjvrsRSpokJ4qL++luAq
HmoghEBeiNuCq6B9SuQeNF2/+mNFiE/hZagjJdCsLOjLksqYM42w9aboZBvFNCB9F+2lUrUmll5j
9goSzjljle5uhlCUlOJyO/yttFHlu0+XnP3TcvBVvqQU79V0vyImSuccMlTNDiyjs+a11QIEZIK/
D1CctYPkdJY/voDFbsPDxvtosGK7u9+X9eN+8aR0v6GyEcaD+yE/oG42ppc7Kumm2zlZSVV16Wvi
XOXR67KZF1zNhSMzbbFg4mSR+d0njyjkEqwjFYIFyyyuckFyykZU+M4xpFth1bjJUzKRgHKTcgsl
JIa6C942g+X/vQ90xzGy72/1uWt0NcCHXiIzcS4hua+fAFi+3bzALFlqCvz33HaOoLzSnlZVPZY+
KOEw09A4oKwzFmPsO1r614nCAnM/NOqicsZWeT35u07IdvGp9H19o6hTjfJKApSkzYPZpZgXY7GR
DmzMrK0ch37N24rNk3Y+pJTBDSzEQ+nd8vfszBeZIpk+vjDm/3Ae70ZLmJ8EOQULo2+WTaGkkHDf
k1pKAEXHwRrKyayczd2gHxz2Y4OC873vVRxChqAnBzTY2FWhWibjAGcivcpayRjcfE7NX967Wqs3
X45qzhW2zncsD2NC8flFsnBFDRPUPtjslS6dV90/rfFJHfBU60TXHFGd9WLiDLZ3010HMLSPskq/
4Dl4WvRKCWPXJjGJlBLMQu9K8yH5BTxC3ty38Fizonba5qbdy5qYxjwQmERV0YMZ0BFWAlcaUooj
O7B4cAJH8lAsJ7fynQ1R/WWJkcPDb/I5KcDdZjLr4+F6CqpwYW61Z14YeR/WqoEPqQoHm+Fqy5Mh
blkrajDlkO0/MAF5/I0lX1kO9p+3BFUObXgeIKaurI/PPx/p+JtIuQ3C7sz6Dxi8nhmmrAD0jL2m
UGLAsg6FsfQsx8vnSMH/g53DdXlAAgGLq4sOvQhIRSEENhlKvmEdbmlIpFkMBQotnChXZn747fC4
a44GVjRn7sv5cnRlpSxYbxIKeHZqN6sOTOZKaIq0kdNf4QebPeBwmKaIZPHpIaWZHo6rgYZIMAWt
g8CZ6h1hLCxIqxGpNyueOp/R6v6H58ZRTffSvHiAwaztTRyt3GSIiCPEhFu9AXRJwC11418m2wk9
sLAw29aJAS2k92+jRoTeTZ+C5qkH+63FrBe3GFjDyx5Hwm4fOYoFak4sxbwdZRE7WuPrEPcTL2bT
Fws4IlmDYBrZUH9tx1KxvDEw+dOA4fdj6awjH5KRn9qx5wjJyTOpj/1tg1xpVKno2XZG/nvqzn0L
5XZq89laCOSlTwUARbEnd7pBQ+s3qUCZ2n9j/Hpi1ozwqs1AHJCqMN2rW2Ctbgxw++zmJ47e4qWK
cwDQTqFLXa7Gq4uok+0pQm0rF0Y5JNhe5Gg8k4hQf24Pl/i6+x5oVLHgdDHPCUQSXZni6zFv048R
79ifnyuXEEdvWj/OTEknTUidXlMEm394nJET5LKcmjgfiFlzIw4enRXT6jCU/T1qDWWm7Z+uR1RN
j7CHIHMoHv0PrpU+wN2/cU4VD0VdxnkY9EN3FN90yz6SBQeCVMTx8ncJLIOIJl7D9CkIZWx3mDHi
8Y47CshUnGXNUFp4/S+23Wre1R+S979VbHuiKbJ5PmGQnAS4V0TcihRw/eXPrFyb2k0nz5i5v6Dn
r2QNbzaaHYHuadWkfzBVYVETdFIJxxx10RbtXRIXHcP98kO2Ori/gWsuHMuX2ccdjz34EjeTZdE9
O5y6M7qpBQkTsIaIvRq1AjCpGwAtQAVV0/1fBGdInKT7wbyQz/Ovdvugy2PTzbuw3bWFkjCj2JSL
wIcJKEuUX/JJMqeWWgL2Ap0vkw1+x8Ggk4IDPvEE1wwsfBihBOthjVy953d/19YR6I4c3dZywEC5
k2Lfj9ceDQbvlkHXm+n2RP+rB+VkNo71g+7Ohsv6cvmcPcG8DqYHJzv6D6huD7GSjGzyZCWFDBZJ
L6F+M/DsrQ6nCZz/CysJ8sMxsFCXPrz+CJGKhvt2kvWBNqKWUGlqo0Ux5Lc8aSOu+1pdECgpc12C
wz7eOOuHVrwD074lduVMqn5Eq2vt8tEUar7PI0rNN1qlyrDJObQch+VelbIaT5gqJCgXUvG5Vb6l
5XSGEYK7MdPCN6DoVT7K4gfZNheu+lkHQdRTzoMVtf+hBUlRytS4Y+fM2X/mzmm3xf8Ca8qQLb7M
NzQES0vHEJIAXMEBYMmt3rlAgOI3baY+jvYw6WpP9/4eRUSUJ3murjf1+jgaYX9OHxn+g1dWhKbg
Ok7UgBua4TqcZuL+GXBhSxBaYOGVQqyke2p0kZWx4Wh+KGHyN4g0COEg9JGH3KZh6Tv/eFKcUEHL
DDWo0wEQ2Ty37mtdYUqP9RVyvFYkv3AihNZUr7RnkfUv+5cL9xTmnJM8D0xqfDGg8GZ8elWIXAeC
65YDV8NZU1+Rb5GCVxNh/FN7KRW4MHaQdl35vD6tfvYwZ9jCaaSK8HkuQOtal4EsFg1qSMCXw/lF
XszNhuW5duADnt604BZQKhP0bdXgHpGlc5OYurTJsigoPcOXTjzpmpwXhVJ9qg99Nf540VFxUqPR
kVQIWPicMk22ALPoW+3WG8vJKOqlJOHQ8lZI21df9KwJcHpA4FimUjYrLG8ymQB4IeTq7dBHWJjL
ZwJGu1r/V39aoYf/KQ7NoIxLHn72RVrrumijzC+4VYV3kF+V6NY1RFgv+o3TGoHF5gUkuB0c68rd
W3/61sXfWmORrnSWekRp3ulvtpMkeqJRaUeqQyQGQRgRYtUykq/YUugEXsxtX0AZESzbpIv0PGSM
1S4/jg5szH+7LLMGieKQZJHy7f2ov8+vo83r7Kjg5ywE8xub1NJ179F0L4JBIkROX1o0Xu83eXRd
P79fwBt0LcbyWAx4j4QZlL6MNFwHP5rwtpPsV65TnAtq9xe3+XWyWrotAErFNr0LumfZ5Dc93zg5
DcDr0X+vcSwYENkCPhefrSwqzVTrHir1bqFanXegqYgO5dmejT6gKL0kLzSfKsONiJwxvnQpzYAR
6p4eoGWQGlMBH1T3/CRgg0+llr52lj3u1jyJW9+iwX0yNHtayrI45dRKR+mtABpFO92e/IgZZKL9
7+QZn2GjqlqhZGKaRWYQsD+1ETLsSitxWtZRmlmBcJLQ967Z0BbeDBJ29Hh1DpHakE4ElQRWDFIO
xhGsE7rOmRFR8jz3wqhQj1GcjFM9WM2v7gm6dGU0UyJlDYjmX/MwWivzxwiUl1ggeQiCYECAgEFG
H09humenW00uZbGdv9MdB0N2bHvX2Wz5BXLPq1XMnQ6o4JSZv3ToDg3PKGK35U7bXuNUWie7h/ew
wc4vCYksQxVtc2MOtjDxCyWRrkfGxrS+oi8TNXN1VnZJ+GKNVK/4HRXHUNnXOMRmUI10Q4av9Qon
DAiUBmg53DroSM7WH4PqSxWW0X4sRv+PVcjA8q6751WLFQ4GePP85ybUtAQWee3BQii1eYoD1sip
wRJ/TZTTx+fvF9OWdYhLoxLmrt0jBt/PtxqzoLDnsiHj5ubj1osJ26bOpJJtwHrumq7KF3Vkx0kr
k7cNiDaVcnMPm+bxFPche7tBTZjYtuwmrmzMTenmyqoVYMPRqCcYVRoHPr278vKsEa+2uhLtf2QH
LnLzeUyq8M3iQwYz6XkoIeKXYBgB+c5B6Tw+NrjsHqOelYiCYMR8sXaTGqGet9PwUA1cUeV90seU
/qOyryzEIkQmCdhGU5s1vLx0CqzC4kWEhMIGkO7MJTn8kgBXnsjg/+YxklBud8H7uPM7V5KR3o7+
w+8fedQGzimzi31oqgdmqgavT7x+kE6G6l4fYcQ0zbXIv8UdiINXkzHfdEBpqqoRyumgv3SI+qDa
C197f6OpLkQDAm8OPxePT3JydRWAbfnfoESOpLiz/p1oi4k46NLi8JNkFiWvh2nyohQLPUgyOr5i
Ss27eFEeF6VcJjc60Fxn9YISFvRLKIY3UDPh4xH5iIGOz/BN/pNnVqPqQ/4Q+fw9FZkC3Jj8yDgH
LdtTjhWRXxKRuPijVzeMbI/Z6rFRg5i6AZ3trJzD1aUS7SAgLHTEYIAUO69nUfl96GP3BrmKYxsF
U1oOMwVPORdLF0eBQ3P/en8gCa2wpUmoZUEzP1ULAzvfgCE8C8sR63Yks80NeFWT5GltoTyHKaZh
VbbcBl256Aqar57prCcY03MaRlzjEG4wCM/LrVI2mI/EAq1eG3yyFT0Myk+FZ20iKHjHDBoRuf4k
3gajPb5LMYSKtcLWbKxnHgxsmGIJEMuSuqppOnR0Iq8eY+5B3bU9cEA2g2OkRuOxyeRYN2CrGH+u
DmgIsHUWdKiP3f85pWVVWx588FlWCJtTKEeAdch6y9o2fvSFkRbHMr5aPPPuwdCcLb5BZXlY/OFC
F0yT1Mp68zOVYrxslPZLMi3RCy2aPfkm7HK69WMcYkGX5ywS3tZlnU7ftAbtZEz1Tivwum+rpaJu
jc22pIC354faIhNRwLTlVzoisp35VtaMaN2Wose9K3p6XWaWz+YZHXCckL4oTxlNL5kXIsdyRvYP
VHck2OIHZ4wx97N+tpQk4kDfe0RsBRMiGGPLbBUAYJuWtHwmXhndfy82Y5AQjlzDVk8oE0Q/CahZ
IfU1ISBCwHtU4DEg4GaIEx/fzfRX6xZrG6sc+e/FefaUtWhpoQOb6m6oSMzBpI6sI7dCQjNQiMo4
1bMDI2e8gxkL7QjAGk6eJWqKCOaYR78wPnrS3gWosSauqlSHTVfaj7QrSg96zXOQRrqFsr2mlZg/
xTFc3rijhpotU4mSsj5uVV7QWLE9kfPYpktsRACSQ61qmCZ8w1qUaYQ5tC/2vyExKvHWT6r/ACKv
tpi9cXD1StdslvFz1KDGTzGDBKQ9SyjgExmRk3dehAOOZKbTs2HFLXjqb3uc2qHjK637jNUs0guT
k8tMQgEcDo9877DKFlRrCbYQtV/ZL4jVXk/JGGWo8iQf0bQGxMd1AxqHT8JzNSKvgzkHDOPbuqFk
W8uroCCYU5L5gDsDnpWMhUmgX22Enh5JZwi0I7nhBXFFcO1x4e6TTQTVWLIoJpxL0T8OFRpdHCLl
sS1MXfiiCcBORqYmflmW9II5sqqGnRAKpfgFwA1B2lZwm0Ea6oJx5UY2U/rGdCTDGSQxVLCu4CmT
CwvlQItcZPpjHk8s3k2+zHGNZOhBmstlkUSujdj/d+CO1zgewQDTKQz8tyQxurkvHbRauPNFon6D
liklsJT/SDeC8z+fUHGo/t1bLg3jYdE+CRwNo3YbLZJrI7vLiOtEt1TP7fIK1J90yAuRSOv8dnQd
i54607tf54bm8aVHZmGNM7K/vhC0c+YBojJ1hr2R2rJjZVjiMPnns34G4UBT8B1XE5xbFWSzCgVJ
97EKf40ooTK1q04Y+vct82zhCToeiLzSbA//MvcUn+MD/7UDwqIIlYP/UPiSjMVBngN40+MbKP62
VdOME/Igk/rD2EywZSc8CbKHn/72z2ygsjJ44c3hBdIFdCx+W/y8zvHrg11B4hzzOFq2wRbYL+p0
u/WRzOfcFvnq2gPeZXQGxTJx1SXc9RB4Q/zdGvRRJuVycWhVrVMdtSTqVdwOgoZJmwORLBlBeQK0
XhXMdi1ZwHDTpF2RJVwtVqeX5Kt9aX6NQ9hHbIlHKK6Lr3YD9mX96ObyXVB4Ue8TdyZ0PNNxAktK
BKzIXLho8U4ltA959l1xa8L32yYBLojcTjMgnYFeVDHMW6NJmwiWs+29fRHf9cW+yPQ7mDtM9RwB
nhzt2WKIL+3AHx7a2TB6se9yGKRZW8I2VdZy3nbX/kNbbLOXhaDnvbOJCMJF8j2v5qGBwLaZaScb
UknXFvk+3tk7dqKo4D0KrtuvZVeJIdDytscoy8mW13vFeX23VymN71nLkQYXOA7+W+Ky954sGgCo
lICUBtqNhvgVaNK1kVXC1yDKDS+tBuITvvgiHRc6PPLpUF+F4W6UU58hOEdUX/lRoYg9AQKU5bXx
QSQ3VC/kg8kg6Tu1pVOjCZFd9jpMAC8vKuRzca8KEbUoKynIBh+yQBjlZeNYtcUxCM3be6a8R7Xu
b0nTGh3Qn+AhytwdFb6RrkAK48ud2oRZBnBB8Z8pGBI7ukQkl3Qd4VadGg+0AqAl22U4/XUab8hU
Q4kn+fdOqnqtPGA/k9sovq/VN70hsmGH550nXrFtavL5t84jKXiVdhyLuwGrWp2I3Uj5RxHBXOgb
21s4sf0RfycLtf/gf/Jqqow7CCNIF9kfWvYTyTGcuiMD1yTetbJUl3PKVt8k+VR6h1UfAQeFSc5e
ERTUnJcksTQXR8b/+Vd8+WkK02bQzee9ph7ZsqJc6qDp0DgJXWHYBjNFejRwsisNnYk3oLblen+x
1hTlR+/Vj/1+WFVCl+EkDV4aiBjvoFXqlpb5NAe9FWQkSU86FPSVRFLSsOKRPV79g2DBXf4B4MCX
CpIU1HA+vanYZ3ka57Kpwp8XofW5/NqgsnfDcJlwjfG4m+/l9AIHYO9z2eNhuA0i86Y+EoWSNE0U
cgc3SuSm99mo/SX6CCS5cL78PKmov88/TzUYk3lvvaqMZa7AN+/Dp5G6TklQ+1HY87fiMmSGajS/
MTT6qJpjdPVkal3tCjhXAZAKxaWyAOWScNu1Kpvx55+Uy1SlwzJ8YrIU4K1N7Bq4hUxN+AvKDZSg
x1xIQ+Q244HBpIoGIxZu+Rx9FyK6pke3lH+f7j2N+Pxi5Q9lX58Za/9a6IjQAZVpCm2ISxWgrni9
oJHCe/DgVvKJD8aaTXsmIUa9xtbs/IoVWwDab+5gwWdnHJyEfk7tpytHJ7aQr/PiyAMd0C0eZ8bv
Hj3f4wODKbUHdn72jPC7zM/8TeYlKCIUgXoAp80SaFkVeqLrOrLGuvTF2PveNDnJsS/zAFkKSA+7
dl/JV6UWb6CHPglEbZfnWuM54i4JYk6Wq8O/ZX0u/eQVLD0uvTxkONksh3KCj8SLel9U17YVG+hV
xALfZBsJeT9IoxpAHobSw167BOgT+dCQquezMrHQPB9XtnNXGh92kwpIGSv+C1/pIdhW8NbzKBHx
Mzeq2SlgcnLebDVdwY9DUGtro3VhmapILfpitsWBlD8Ltlz7ERWjNj7f7OlpeLhyPWKIpkqvMJ0Y
7EfFACKgiIutbMDe53OCiP2BaKhpP/ErjUlyi92Wf/lE2xny/O0FbABlWAB3fsJSTSPxJZF//iE8
ZP1TWeye3n2Z34gPQiNUA453euLnZR862bcb09GnlS/G7W+7fNLMnuSzGzyMz+2i0kg/+ouv1f0E
WVt+x8ppERE8u+J2yLioUmpihKhJdQvb7XsfiuZWFIxTy8VjwNW9GdGqmPBW+zYIJrdxhqwCKgf4
dnCFTDYXEi43lWa/2lPJE0izCyIxKfMBAK496IcIIkAsOSonh3A/AoqDescOCjYwi6nzY51Tyamf
3c5H7ZLev8ktPeTZ6n5XH8OQvj4MLdHcSDWlCugpaZUF3fPyC2aAOlrd5Sks+/GiATLM0PhhOge8
otcdIlkg2bFg0Kzyf8pAcXMwzmOKCzwgSXRpn9k/O8qhvjV9FSi4S1Uhx5LW6zwdDLyNWjaoXvPV
Lfb1t3FQMRe6/TX3aAvXpPAd7gkICyrC63tiCBbCN/aANeRwpxahXJef3K+/fmnPrBNCJM/P4Wkg
WSENKf3XND2E5yCsKF44H0dzFmqpJhXoA+AOuDfcOjYOPWfU+DSt+yQ5v81PR5xgeyZg3kBkQQS4
tv2luMhnjyaJReQ2wAMSMdkrYFiU+CNj05KamjDeXaBR6khPTxooQzFU5W2C492I9Xgyucu+E+4+
g3VI2HdXex7RAtAAv5Ly1a1lo8jdpc8fYnK1d5eB+E9IwqmotM2BuC0h4PCGUtsyMKISfETuzT9S
Cy6e9LKKmM9R65yhp731MiUNzZhqIp5TA0on3ncrxwuif6ePh250Hb7hi6tJRkS7EsvJ55kv04Mr
hmZKTHyZhg44FrhGvGoY9YjIN7Yhw0p5ALP2hPJyUNM5daM4mo5qnj8XR8XOzes6tyFK6MWyI/hJ
VgcACMyXJmGLX1uGJScP8HfTKzTTfkJ8W8Ep9Bsmrj2m9z+Y37t12i0xBfpnYkbTTQnzqnh2J/Jt
8S4Ajt4fAC3MbbargIldsK303jHRtKRG6bSeSEqCh7AXAh3XOisUfiw6hxcgbqQnOgON8RQ1FeMx
BzpxZmTqMTDzGMtEAJ2EnCCudevdXZ3NyG13o+zDlzbtKokVWPp4mTqCCiqBtUcga9uPi1tlyBXH
rdbFHwbhcUb2h/qSeq0JtY7z6Mx9ovYMpyeF7fS1M+gVUl17XDMUo1ip+IGLGOHz/ClEBnURZt0p
ADwmt+ojdbBcr2pKyF5ROn7pyBiht6L6iB1dIx3H3hZWU6k9W56kTe+PIi+wGBCjNMovnjV8kMtK
P9eL6xbZLo9fJtHFl5v1NM/ttzhtabHIex4D1s0O5bXMSRmP9T9vxlRrRpc7JpGLDpC9D1WQXP2I
k3yK4wlnNhuxVZiJr+CfTkP0p1nKyw9xZdKDzepGam7GEPMB/+K1R5cYvmdKEbUbG/uGQUIBuOLO
aTJp3VOBwXbWmte9wUaD9Xf1hOUMQm0Ega6OpRNUN6DcZdKAwvukPis8z1ltOCfyAdAbULZSqRha
p0VtInQ72GlzHN34QMmfBAPZKX0hHGpKi3MjP4gcV3vSHpJjuh6TUSjp67xRtKFtez/eKyEGJeCz
3MngG9kDMRe4HYClO4f0bLC4BW/T7iz+4NLXSBh/s5eXWh+uzfgGr6EaCshY01o3P5pJBFaZVzak
wWsuyRmN8mvvSF78tmA7cL7bN7Qp938YA5Q4TWNmXLB9eb/OFrD5Zh30tG7sClQ8+2j6LUikrJt8
kmY52laI5UAttpENuaFZLkY4Gd98DEOmkUc7diaFjvtyEFLKNQ0Y+Bpt1/ARW3Ez7k0u6aQY7Iwv
dMIqXFhiJR8k4CRsBD2BmJxbQUtslaxLL/NGSgTFlFDMJsdeNIWPiZSZodctlyn83hFBHp3KJqe9
jbWjuR6dDwQtSK0QcCMFtjFBroku5JgLmQ68gDP6P8ZT+x606xMiaw3Udo04xLcIGUpp53r8yEFe
LJDU7LtOX7ztma/+vfC4zASDFgSozPWKDo7OiCaESiQb3+KyCeZFWn0Vy2AdZtHgxy+ZorInD1xI
gMtBmHQDJwAeU96KYKxnfRNuJM2vY54ZzeRXO+Zd9S18b7jcV/QKfnfr+HkdLOVLyIjEH7MhVHZU
DGhhrlUgGFtBg4+hI3PRPzEeRnWyQsmvcSLx/UBDrN4iyU/27kBd/VagE2ZtThkAUPWnLSiuwJ0m
x4D8l7ih9PE+agQ9cbC1OVjuWX1Ws1ujZUB56XilgZfmfDS4vbyj1VOclXgSjPPxuDJ8/W+Kyx7r
L9F0m7TVji89jXX7R6kAS/lponGsjk73tJF30VGz+3cQ48u665FbR6K9Eu4jcRON9SvCCOfc25KB
4ZJgjlES9ZPdzG4SHEMBIBfbBQs4GKcasiEdq7MebWs7z8MFVq9JeLGJd/n0VhChtTn3eLiTaiBH
bJQN1clEjbfaxjfUcm6tzA3A91yqa8PsFVRRgdqMS7dj3KMdD/cU07rEWYNWSWtLmoCFRQpHhs5X
QgNSeJHIzxMnSVUt6A3vFw6RPrw9V77ufQlJeF6zlTfBAhcUJokJksW2T7wrXUiGInz3du5Ol+8k
Yy43VBXSEkdyEI+B+Jy1a9s5CATiIreDzo/TnSlgvaCk278KdNdgA2EeKVpIl9iMgndOKc2xSH11
dEzN0gazVY72ywsUsqk0ifJjVfGXDWQlYY9RKiIHxLuYzSR6MhN5U2+p0zJ0sp77TS7TwugPl9kP
3KsmsjdO1Y9iiWyqo75+C0eha+LEk+fKwAKkIxDJITQRtJxCrculDty1/YrkINQ32bZkizc4quv/
eW3RD3NjHtj0ayErpTxBRAdmb4xWe58mkir723vD3hsTitCiWVrwnPxM+jinkzdSZ7abIGATmC/6
CLZrUi8vijGvq7Fo/YBx1tFB9rve8MtpGd8xOddiQac+S+mxg89TlOLQORlrNvvYUa17rvD5KzHy
6+WiDI9GRZMBQaHObJfIuRhTdOmCEDRzUiSX6yGn2yq98PVFVGif8hZIXNac2WyFY509MwbAhQe7
R8fSvRWtWe+D5qtMVZZGk9LDFk0YO67DS9N5VAuyOQEOm1uZd41hK8TiCFvbxCn7NPjUbHYt+SpO
wI74cgzzN6mEAXhWWTinRzS9agjCMInx5PO15+iZCJa5KOE669WbvN7+09+idlnqt/KmNGHX4xcY
W3oAb1lI/WWwzJ67VIHnILuzbox3F+dY2ChTeZ5sjDF6/Thvg/VglP2WQNbHu+8SBaKVbuuM9bR/
T/CzvbHViKpX5p/30ZRockAA33C0x7YL68zTSw1SrexzslmQ1TDlq5NJVf/TovZDjlbfUjVUlCv7
Qb83r69n53vuxBAtfhoLpT0sr6Dw7z3Pn3yZB/dnUHxdwi+r4bNPj4RwIycy963qrFt4OJC+0Bu1
19b2ELWpPOx+ulvRGKpZFLmmf6sBlYQq8/m3iQTchaKqM7b81YiGMkeqwm/JcQrhsbjYna9GZ3r/
Oxf5qDPCeb5MwxIbqKrdjF2UymxTjdHZXEg8M2ylLZcXcelydePEopTs2vW2HxB8spPPYVO7zy8A
If9/cDURcjyAqrskBF+I54x09eThpKOJ9Wo2F4X8mc/j0n0q7E37ivQb1Rhpa2tEGaBw2ris/9Pc
PAoB0xwCseJzTxrY9qWdXU65cwzfeQDe4aS8igxIDX4cDCDp/2N+yjoXMsoHzjLAZWf1rhPVgB5n
YVsH//dOpbLSLOLLWbj1Qq+OMPyOsjRkMeNA7hYdLFuGv9dyzwZJMP5SzlokM6i9QoYbLApfLNCb
e9x1Cov31Wq3CpaNChJdWmkI+T5u99ezFXiQff/7rfP1R+TDeD1V5/ervIgrQR/UhLH+UDmKMelY
QK55U9ehdhmFCjS6HGRb663440OfZSD8R0wPdGEDbCsGOaU1EVX0NWWGbOXRbhhEo/tgzlNSin8e
qo1xs4DvmTPAf47xURkvtc2qDpnpYecILjMEbF6nZU6uu82e/mJAKGvFEfOW0fGqRGmhBrnK1wlx
9+8HA4MhSCiJsiL0SXdDfL9oLI8ziK/X5+a45yq6Zu00F913Z/05M/Tm1C07KIdXIh17/DRc8scc
9Tqk0qjOsKgBKN4XpL5haOwVom1j1Rcso5VN54BmFVsX5s2QIG9Mgn0utuiRGrjxqMEZEMzNt2vl
T09ytiPw2EXS+v8kzX/IgCZEXTmGismsurBjYAljlNZq0Yy853yEOZQbUvEmOZedY8IhZJLzYWiO
YRbLv2s28eCDb2rvHLLAsbc1HRH2G9cKIV9YgEDsH00zjHOpFoL/8bRDj7kSQG9C2Fk13ZWWdCfq
Io+q5QidfakvJycE2y62xCuEEzHN4H116CVXfDC7pUWXAbT8ZwF/zKRgNv7azCljemP9I7hVzplh
L8SXUstBKJOaAPdq3CXbz0LU+M9KCmEYiVa+NGB0d/E7xQorW/nPAHredZ14YRTOwIj9ive/WsA2
bhL/NTbbUUgA539uH3UNQ584a+NtX/UJHLIRgYu2EPBmmSUJ5Tf4voR9A66tU3x1AuTDDDVtFLlS
mWchr0Azg4E2AD0Btqsg6jQFyfCN1nu8FiY8lkI/0698g2yH2C0+eXmm1Ms87UtUFPXJn9XY8URP
UOmE12zYszcIOeJIVyu4RoxFzq+AWgbZqiqixStd1oRT1aczMGeu/zXYCITtf4P2dDAOS/cRsLLM
yXWjAch3WFrzVVAqdZV74+JP78AUsFONc19mTyGU2wF4S1PECNLa4oZR8/Rpb+L2V9CNqo+Zp8MJ
5ZvUBpTnye5zmq5+zMTAhNfOcTtU0rZK8KgZ0B8wY8VpJd52SuVsbX2Hg/qHb2Xvah20P6SCiCBR
RDtBDNhwzaP3alGJM5mLJXPh61B/mKQWksx57aFT3SWcWw9g7ENeRa1rT4NGm8YVlvIkxVETg+CX
NNn+yTUp09mIX5Mjp4TNVA6AfTfzcAYO7VexlZgm8LrF30cAW7y4amIAOYiwRxN4R3R8ONeGlGT0
T6Hdt6QVCUp0FFvJJUiyLf3ggxzPl2HwNixmRnIO2ZZgp+NcgJwuRRNgi2GDekPTlz+VnkQAx59M
C+xeXQ/hBm/40RhJl97Bafge5zxGXA0eBWZ2nHef9mGO9aot7eTeAR86aJvOBkaXT6QE9z7LqPjw
ffdJpAloMJbBCgDoN/hbXm2+bbuCLdFUC4avw7AhXTY68G0I3O9pGJKWMuDAUvUKtqALyYy6tFlf
zaZmdzXYvBTT0Mq+HPlYjRlT4mJkHxGl7c/32lejGaNKHx8wH4sJBsCpTOp2RW4hvMCCjwplCpEJ
kNOJ0Voj/CcHs8aCPdzoOkzl18J+4qYp9YQWbJzmP6IzTY+XjLJTPqGYeHGtQktK+owJ0nrlvbDV
dTavd/bliWsXm/GzH+VEptBSV0K4z5aMxU+DEGl9dHkKANaxd1PXsNHcBD2BiSpMM04Zibx158VR
hfAPBDVMHHPsdcQyfRCgqKqbD9DPkFQySlHHoOHg077w/sBQrU6jktufa2yirk9JKNL3R7yU29Im
qrzk0gqkRrRF0sj81IF9HONoAJXJDm7Q3cEzAVYdX5Pm3h9Q7XqAdWT1sqq+rgGjjhq+3pL+nE4l
VIVPJ4IuUL/eUhEQqMuewVzP4VjBrQorR/DR0G15k44OHktqQxBxsUk9WaOoS2fko4Jubpad832d
XudmZ8psGGKUrr4bp13fZmo6w3Ack68MX/P1FoHajt83ejcPnRQGzl+8I3FWf8VcTAeevXUFQPEm
UzlCktA26fAvKTkLsiVcaju6EdleQQdDPnxoAwji4pl+Xou3dCUYEqeZqcYS0i1JUs0jDRo9C4M4
PBOQs+7r8uIOftaYFIDjiN1if+cNqBpYDGkRnPPG/7aOjip9LS303yJvZ4bMobbVHs2gZFtEwc5X
Xjc56MuUwtK6JEyMPNH6mmS3fbB+zmqoDEFIqm5a5odZonz3v3bvtYp5SeRWeYKWtuOIDKJjXMLP
3/hySouPqfaPv5UzUerAxzMXffwEQxyq/qgUTVeiaxHHMbMktChBAwiVt+v8DyR5rSMB3vFjqJNh
8UAbt61Jw5eQG+fzPvCIpLjXlAp5FN6jikTrDHYpBDgrYT/y4sfAukA6TKO/Lz787qQ6rbVnHsIy
xebTMpCb1+AFf6DQqRLeACc/HUzr37bhH6s6T0kldtk3p5c0a8dTcmIlrBKCta1+crUTOX09VXJF
av3M7jCp+A/rpH+qL9AV3GavVj84kPHrfCG5T/6KZ1uxZyIQhpADgGwvaDM6Je6nCoGetKK99co5
JcVJER4dHgjPkB12sMGJedAV+yB+6kz6QykY2AXL2HQ/B1QKLGwqBHXoR1PJAwV0mrx8eTYZkgqI
4P/ecE43R5iqFzMtmlXr3RJmxnvhcVmJVgkLd6IotCo40HEjKrUwlpm4xGwlWk8U6oWZ82QqnmWu
68nLGunyfftosDpxIw4AqrJQdL5JNtWMh3TpGSqq7Cp5V95ZByhJKFcw7sjHsNbbHkgJHUUrxcNO
y/8hiA1b0Ptnaj1YDVJnTEcy7fHcSSROctVQ0fan+YC3eEzp4wU6heagvGy2J0Aru1eTp/Tibw0C
wO+kztj9Tg09p1Kv4NhluxNIttVGwXlK0XSabxDieYMeqcjtto8KfSH4eHO2licwyq4Sa+0fCw8r
bc+2emycKZzAJHddndRw3qBTlh7SQ9MwNlQ+KJt2jzoXPlfcHanpmK1s2ll5cEgycpEY10HotcGH
8Pp5UWnQZ7tbc4G1uMcF+fTW3aFOPRPkiHW3wbd1VPkFd5+l48yQ06e1JgbX55iNtrhu1qdkxqUC
2Tk+XrPgDBRj16nyXftAqFUUkzRrQwEpZN/863d8myPz+w85dlr4LY0IdOczINHA4Q4+SYEK0GsZ
22UNm2f3mfvzSqRqj2XhwuK3VdgyaI9iTqLlqtYQ6XdMHPhrQ/TCnkGixAVaD9jPH9XOQo24k79C
CAJG74mWfzR6i+jNJsfVh61FXs6IxgB7Rztx8NP4nuliZThF0b4T5j5NE/j/mt+mIPUZAR2RTv6x
LsDrsiu3traaXe280LE56z0km9COGEqMMTCJ/3bVRRYehvg8BDjlEqriEy6UdxBMgEo6VwEMNLiv
R6maNKF6COtCAUUv1ec4xRsqyajzBCFslTJ7nOHeEBSSudMAkbl0sVHYtFnOBpu/rVqZYEIAyX16
gElk+AAWUvXnKSEsf3xAZ23lqGUudZ708FhacpWrhbsHkIMhcaAAhk3kl6YS2UfokC1hACbnihzV
ADK/f8Q5JmvdrF0SzKOrc5DI1Nx0UrL/X3G74PYEbHSlUflbrAvFuEzuwMx+2WBpS3EopGgNpJoy
3wb+NzAeRobujm8/kVpyvOntolte9fMWvlKpodPlmGi5nDuV368vP5ReYAYV5GEA/xq+O4C8/wuK
4jeM26aFsfIDUCf9ro8isaB+YpOkEikBKbhXPqWrKyoOzWhYlNKJdd7i20lu7KD2pyEfC7AM9f2K
Ni8+k6XnSlXZVpKXlS+zgtOu/teaENK3rZZ9aqQbu5xImzc+bskKNq1cIioaA1L3FggNB7rj1g/H
FWGo9OAmPuEASGSM1CQ+jZglljprW/3hB9cdhCHpeUw3KZVYbRa9N6x1uuEupjYwVFCFQVmV6MUP
HjZeTP3/G7aShshPyz9cKjDHZgTzYEFRh/yVhAqiUyaMYeHsMtVBXsbSqEx6d8CzCKWv5Bqz/yZy
61dY9mfDnqtSZQk5XdF6TEHYaePKqS7VsLuPQVN8DHvYTK35SOYuSYSB0G3UqmjyQ2YuCbFLECtC
L8URtgybx4NWaeHw+nCkQq32JNKzS8EyDDkxjT2MoXI8gJaNOYSZ7mZKTNJCKXSDEPFu7USKCYYM
E141xpz2vALytX0suSNO8FRQALAEoEOgce1ki+quUZc0hu9vRY0Pmn9GdWXaYJ4emMeS44kz9+DY
Mbiy++zxnRvmLLhnbB+selTYVrfgbZeKolTLHwI/oDkX74XC3OUskDBVBRqHQfqzRJAG/PrT02o0
6SJdgmgAce9PsACYxUa31PfPYlnTS2WSvV+e+K911CIwlWdxd7E/HId6r/RqnxTFJ/IGwTCh8e7C
A4u4jRl6khlgZxyi6Ig+qlSO5vY+qnC7GjnokjBYei5cQPGE9kGWUmblveGNq7ISSf3T/V05wx0s
bqJlUnZSf5g0DjWpd+XG6AUaCuXAXSbsZgtGQHAY8I6oQB9MZBYITDtx0UDQGUHI0xyMwK76KndU
ysQVL8E0Vp57ZZQpuuPGOTHQtTumL8kcwfyvVlwKhrdXS6fVYue3Yh/MLjVGKTUTen8g6Or9FO54
phWYZmEejiU9W4tF7N4sV2X5wZOEGNI92oTs3k8GTFMvWOw36J8VbOSfGhdHniOogLCKi9VHxvV0
83NHAbStonhzZmK+vMaxBIEobJ/gJAxCB1cNCtq5iWX9rTxDgICkRiUxbBBkfbF4tHwbvamgsSpB
e8AFgAVruWxAvLvBnx9QNJ0OEWS334thOEUG+g7cLXGvIvENN5lQKOfr1kC93MaPdPqziaO+PC3k
18NLZ/dHtVbJ1rMoarFBbMDkDaRWj8vcxWPDQ6zKteXb4RbQG7RWGhmlEWAO1xAwSTYQP94+VkIy
783dQ+W21NFHXeXtsSPjM2sy/XsLDS6eldlwinxvja3GU+R14ISx91T0hPHf3mdjuKhyxSf/ydwe
ABRuy6ZBoL2p58IHLRjl6eo0++Yvma4ae4PtdaGgQAac0R4yp0rWpKWXAqoyb4JRCedw5E2CY2Dz
9Vi4urJaUKORsE05T5ga5/bd+QX0pv//Y+NwGl3x4dmTLy/11QXQmSzE3ErZWwb5Rcq+6cSVNjhn
eSPs0dzy8nhIzncVXtF+/AKubBvg2l0K8Y8rHE5CcFAFLjEK1vI1dsP6rVvqiZBeDS0/ZVMKaf9v
ny0T6/l2hQi3p8omnyLxWmocDtumQVVKfQsMaZ3AsFtbK5Mwcjwxq0xol/3gEIBROsFl2dSoeisf
O4gX7Dt/zeXmTK63UxFq6VCA1XPWVYserGUZj0RvzuEJsLL5utCFAWQYtpQld7x18eHz5+3QOqtu
keYXDN/Gxzq8VLsHf32hd2f1qt4LKGP4GoW/rujMAI2sw38MEQPTW1raybTTAfEgJT/V+n0hgDqS
qEk3hZLXIoSzTR4BqsXDW6DzpNlofzOd1M5EC13lDMA66hDpAxibAX9aIWlZC957XkFV+/P3b8Do
SSsKENa/RQJawqF0KiXz9xVTm00Y6ZDog9pLlBGWczCQZsJA39R3JiD8nu7cyJKVNMXdoK30H398
W8eZK2OuYRUJeinCD423RfXgmo+sZ6YgvKcLMKXZpgWPcnwpc+framrPMrnLDxjx68THgyXEZAf9
uTK287wHckcqH4jfdqqTA1TWSA8lyO5tTkVX7pEhsX0/XBKLmSJSoLJanLBE779dZ50SxZWyjP0o
L/X3w/NR9Zu8BdArTwCR/a8UWu4JeQ0m0LYreIdX8VK58fQIq57nvL9k/hkTdpZ5/q4VZi72qlmS
M6uVRTWGebdnT+rNpxQk/fpkFQVkp4MccwQtJOIQ9pW//P7c/UW/rq7d/bt5OJ7z4TwyKCdqtCqr
1848ck7822vVMEZHiU92E7snsX7uq8fp47gX0Or6QYzUqE3IiQNPa9aG41wr6VgCc/4ZqFjPEK2h
KyeGYDe3yShTD51ZwxKWxbxXtwCfBnAffT5ImXDj6rQ20NmHOh9NcBHEhFtOitfYDJvVGcMvvLy7
N8cwR8Bp5fKY/+1Dpwisg8rTaMzhjIO7iizQ1WklfOWl5BF7xVUBpkLrKC/zkJ86LmB9Ex9h52uS
N0RXSnHRV+B1cJvFSEmvoL5TsdNCT19zi+gBdj3+c3AQ4KcUnx3TFPHYibdl8RQ3sXs7rxfyqSIL
tSxUC/3ICEBSh/r4vP/D/ya5lhz/ElKG1PjvEPr8+HnzlSepsjbQ1iPfzmr3SUYbB9pkoF9cRImT
WbMr1MjcPgvr3bMRgB2qPVQORP77mxnJBsLQ0YM35V/6Ak6llicnBH4sWJq920vWtzgg4ytbJYFG
RPSO/Xnyje0f3ND/fEbLbeNmcvOX4g0GewgVadmweYHvvz7y+c25RNyALilePPEIJ0+W8giEpaFP
38GaQMs0A4o9FDPwvztR4YG1rKkiXtKJy3wwzJgGeQ5Y65cAqarYBXHbNsIy7wUGcEAwR/rtPyNt
v9iqthk4gAF/odrGX7/gfsFXidTfpCvzmArzHC2S+6jkGNelp/eyP4kkDuewzaqCl/c9pFXKEx7J
NUm7jISU08cobYQp/Mq+i7Squ20mgKLWDuX3fgSl3H7zS0O0UF/9kvS5abZqZn6pjhTKa/sseoz+
iRY19TsqPdmMfJ+0hgWKebJEyTtLaXQa/f1YOrp+X7sl5wrIlka8IUgiiHhSwZNLbVV85fmPwoZY
Z2g20XyH11SLEtuUPaSrh1p3xjNOtQBbhTdp0qkYytvUraRtRdgjOUtehCWc4g6MIgDD+Bz11f/c
HPIkS8LhsPDreAmwrwpdPwwakgFFdW1KuBwNCyGkttbojm5PeT68fPUFmhOjruK8h8kPGRHiSCJB
SYIjOVq+IFDClk9IR4Wm309H0xa7LHR9wyrHHStF3VpmXjeFmdDiubFnvQVJZ0ZvZGsXJ9OU9WSf
EonVWwxJcPnAtPROyxiWnZF5/oDsSFWKDDmgSHfHmzxGnHO2TaIWkJ9kZ7hFrIOYZRgBsMR+XQwb
l7OFvpk86Xx7ryF5DOlnUFAjE6epk0qq1ZlITH2A+djCVR0/R0lpTTNcvqZwRcyh1iibLiqzK54k
z6boKI/DaB3wXY1COZuRZmlnDOG2+Q9CeWxsqTnJXs1eq8mmjuPWl3AEj+DuORGdFeeV6KFFUBHc
F4imRhO/FjQHIXUWfeRzp1WhjVqeZ+sXyo66hT8UgB5Pm8ABE/lKu7EY4eLJYBR7oLIuAqXsOItv
uwIf/n357f7cixYnVQzOfJTRxaWj9GW9dx2eukIsm7p4NZuCHwVuwgQCKicvD5IY5bhPUOkdV/la
eJDUFVSpUqqhbIhsgL4Gj4DUA2559WMqsJHWbBzvV9kthGeCR6B7OorqJ0L6qe/F1tz+wZcLb016
EcJPPwIyhsJhZKbTT5xPqQwAHSfXQ02eT+N9Mj8rSe1djRI5COTotHclaBiNyaj0vAA22PMUwjvy
9rjlE+Zv5RhgD8Bh59oONgQceJtYB+t3x1NkePc1yFoHZEeliVN18/Ig4CrnVa2LDGU3yvTnVZA7
e1ixWVVuXRQ5kEYEy2EAc/j7BWG3iZgT+PnOon5IrGr5MnUoG8cCpYyI2mtm+63SvWa4DIVZyJvM
AlLcBtpQ38zJnucqA7/SWFMfDMQYIKS0tuSNK3dFQau0u8ZMZ6r/tYCcJkw08QzQklwpojnppvii
7Qwsm9RhsL7RFATVXel75fOiog7w1HANs5AHVAE/4caK6O1oN+v1FBxBCIOa1aNvbhrqc5NrPEQ1
BJJbKJ94dvkjqyzkMlGms9yuDamM32sh63T7o4sPhGnYjXvCKIyGP+zt7vBrZuDwXzAICZpQcs2W
DA0LKyy7GnkJAshSQreGIWZv/qVKwYfkLYQDSKCUGiwEsy2Ia7HYF1GMPpbZfjaBdIfD0q0EIL5R
uJp96qfx5NFoZcyu1N1Du9OeDBdeptZXAkfNPek2yOTtvK8I3IOLAl1kLnEbFORFr9kVnPqiF31C
CI7joIZa+63Tp/UlqoV9fIjAoKQgSzOeuFiANGKBxx3WLOe60oWPOjiTD4UDgXf9x1m05nt6NDwe
wn/DMs58CooElQkLGcr9YbKyOZGBxXSMjo4hTeGMLowAtcfFhQXcObo2Xe7T/Ea8CzOIKOICKV8l
oxHR4H+iSNPe0ZIAGDF0X7rul25r+17jCZMK/3wLwqf3SkqezqG2QRZ6JfZIAdc8R545M8mBvx58
Bii2A0y0bMkz1x2u8c98Gob4VNTKnBmi3b82gjTmqdOWQ0ZoHkqUAUEqhQCzvwmJB5ZTMwNwc+8Z
eeJbxRZzE365ipcEqDcDpa4NXFXk8ZmlMEmq9gvFtRLknU/vpjFZh5sgKKDLX46okYEkAqUOOlYr
rl+uFBxkTC4UMkdgAlYzWy8rwv4olC1TGKQKdUX5DhgCel4XIYFG3jPQMSLq+f1NL37kKFvDqepL
6TasU0UQbJgB4/2TcVTys8QKirxPtQSJJeeALeWfWHKXQ3GIELcN9Jp1SmbSnHcnHgDUNp3/l/9z
nLnA9EfPSU7I+qjDCzstP69hv0vGQ9r0z1zOB5+33hH1Bob2QhnInpTFo4FNfaV04tIinRvsU/l7
QYMFsoni9ASb8Siq5iSvUapiGU7sbDmBpjo6+qfTK/QHKM1NFYjmCXuMK6PQIek1nxh7DBUxhcUC
KpAZXAokOjLyqOuE5RVEfM9J6GUyJT5b9r7anXvHx8m565WpIInzR6uJogZ0dd2Ak/HUf9+49/YC
WCZAoaAD1TrOjQ7G4OX3tSQCJUBfs19NWgYEOfsLE2+mw0mOUCMxsTa7zK9y1Yn08Mt5u2VQvo2N
frb1tSAhImAVm/gpGYGzKZuU49fHLtdJDE63XhobSFBZPoa7g9jDNbAm8DZjWk3QuDY838lS73Gs
wO/IGocTIH7+S6eCJ5Ju1gD0/dC/FFFTAvKQM2KgKyC/Qo3KEcCe7znlmbLt9O5SuxVcdDUOJomA
g2rHFvbYE4Dsw/o7/EUOx7ssG2DhojWCBdNco0EnR5u+m1HiD8IuZzT6WEe9FSj/7NvUhdpzFCyg
EdXk6FTOiTXnujdQZ0JtvSRep3sxq2rk/0842yusoN3geusIyXbjoly/MotqSq9JUGtzfOu/oKzI
A13Arjk79CJoHTm6wsw32lTPd9lJQSqX+FNbaHUG2qtSyELwMOwfoMxx0DC9JgrPUOota6gXkQau
+kjfT9JMQNMlzAr1yfS4fXcCSlJmVoBkpNKK73md377fJCq2huWivTo7o2Q3W1yEoeMQkQqb1kiL
xj5RRgF9D9qI3rVS3bNYzu4VAjLyZWCRkbuuHCaafarkveLvhk7ZiGciNkV/C94KPiMa57zlpBqm
LhH+2O9ecxsFQhgIAXmbDEbeouAmIu2DiSJq64yF2CUTadFKGohw9Wv1VNPx45vhU90tzCpbP8H3
08VO+EeM/zdz8AfoLt94O72LQjeNt+Rn5bnQ2kdRabiw1+tSiz4P65FJSjAenp+yV04XMOwaQ9IE
a9LpZm3GB92sUUCAw+bz4khe+m3lI6Alv/YMMKNAOhBVGml9QUWXOSnUSlYJxNvDHdNzkIjhmmyj
a8AD/kZvrJ3CsrvpUQcnpeOFUEFpypkaxas0wWLDntTUM1SPAouD78oMoaAM6YDvZZrT6KSunEtO
28GXvCTLDFBoX6Mi2YvhRVgSbfFSUFYVJvuso+pr3/UxM08y407DY0qLr+PTJZsKtFLhEtxREaKM
hagkBZ350keYYvq4NmWKDz968xo/m+SylXZ9EuMvlRhUAy4Zz2UAE/sGZivQhhXZax9b7aPdc0p4
A/OEKZsYDYnjxonVNUubf27qgiB3ql/SZjQP2UVwZnD2WECclyZv8ZDKnKWoWsbHvvn6Bvud1Krr
TyjmtHYqYSlTsF9xNN4dkgqWdIKNnXga+kwz7hoZkta/sGPAJ8bej4g8hQiYa3fTTO92MpOpuNdn
WLUKnBgvGtz793gfNFRkS/6HkS6mqoLwS8ih0AhYfSXaWtOsO6E8KQi1H/eWXd4b/ZF4jLAKyWRH
25sbYE2/PPY0BufwuTcvk2tqWdx4cqZjV0oMqft863rMs8B+F3IDIhpgxNzG+BqcAFPswuswKu9S
JNL6+5rAtb44W8dTXcRGpjIJEpP6usOzjDmp+fKXfLWxGIOPm+UxSnpNeIKAOVQ/2jX7MdzmA6sv
szM/xyzX/DJMNfrBuzuZfX0cX1U20p4jaruFs8DRkTk+vpTvSvzO9FT/hWLBtMyVbQD8IfvvDBXr
PzVr+KMM3Qnp0mpe4j7ijHmG0bOvpDmRKv7ssCNWr9fKHbl6QJkLaIGyhCu58giUjbmOBc0/AJ+l
J/LKUYth4dHc2J2vdmZ2EU6gp6jLsCWf3W3xJCeQ68DpbAYxRZ31hwzIGG5IRhi3lKIGCOYq79dO
+qlA9YDbgUns7AgnWFZy+5PtdEdeslxA8NHu2nkMsflJ4hLl18WZ0zWI4jwwfWissl71RK95VczR
3IY1lcITEpcEeCFbKSQIALzUMQnqEi7PCoJ/VXvtFWvP4RO9CvIAc90C6Yf7Hsl9c5OI2Bp1poLz
sRD2Bluk6Kb2ln9YFEV84DSLO8pdj7dqp7es6MHoQchS5QUG5sqWs+G/3KHayPA4yVC69KYgcwgx
lly2XdjVveJtbkUSDxVoZ7czB3dT87yNzjI7njNvbmd5CNqj+jBKK6g9IfAOnOzH111hYpnS9g0o
GEeg1D6owlAGh2w//OuB2L+jTSpomfL1qvOt9hU80nEmZgC4rsdOLe1vYCKnXzCrSB4OZASa3heX
HqJ10vSAiTL3Mxne07Q5fmJYeuMfI8xeqv0E5OFcqc54+Ep0iMzzWlR4J0sI1Npb/4Vq/v6UdIJb
u5SvLhrALuiTKG9n4tTXXWjzs6H4KF1fI2KtkJs0wHAnCLcaCWxOn4frj6tr1Kj4csXsBS9a1G/p
EOIUgOL5c2l1EAJIhw4zsnn/SfG/REVnf6niuXE57n0pVzC844ejQ/iyOqwKcDv2vAn9f35MbtmG
JOHON2TxGJ16yZvL9qEm0sIrZYoey02Vi6Gy6/Fo8jvO3+PqLb4zEcVMUCYgeqC2TnOwQytJ2Xd+
T8Bq3ZVvEsPuW6AHkCCEO8UCqz/ELmX1U1cjCzkvmMsLJVCXyqPrrZvKTo8lMBO9MfxhFMFTkogM
PpdtWl3GtQyfixsToZdqwBnAr3jzylpMBa8NQwGu6XiPDZcInWOArlIwpPnz9dEktzTomy3aI7U2
oq53ktRGh30kAnM+AlvuDDKol82ls7nG4uMi9RHqNA1os0eH0jiJuw5hMSGVZ/dVBCLiW+XwDQIP
CZm9wDtDYSSp57HTJ8Naz61xUWIcHMMp14qB9lj4SwYPA2TGNWHgyLsimb1RXNcFFV8T91EM6IAi
kUu9Szb7oC3NdfeK7+AubLB2GmbFOivc34kdylXcjyJc74ofz73L40DGV/Rp99vqGe7WGaMuFoxm
6xTvvAXbXEgltZaX4/PEdf2XzeVCC8QTF9wUa2nWOAkcErNBIVx3DjjRO/NOcDKeTCzHiKSb6NHI
AIpFOa8UISCfMIfb52tHy9lK7fha44mkVA3xZp5eiXD1bZhDpWKs6PWAQqd064c4EC+DMJNlfkcQ
976/ipBKC6aASUQfrz4sY5Eh867IzB/1HwpCGtJoIhXpfjQTmxx5LRKfe50sHbnGGKvPdCccxX/B
C3eMBa9au8O+7EBOv5bhak8DLlzq4B7rIhcWj01m0GJY7i0hpCg755fog1wfqtUz5B1rodWHTk8P
47J2eJGpg4wph58POrL3bL7kNwktCacOKJJqA5EWegUUb1yHj4f/v8/Bas5uTCY4n6o/9D8482WA
GTDAmz+qRi3Wso6GvVk+vLum2Hj8jKW+rxxbqp9+ATtn88p/nx9fJ85FSlUn6zOOApgyqXnS2HDJ
j+wEwdSchxnKj5lIFdJKEYD9hKJaP+6n0QlHh8slzUABINRzH8Oo6wmyLgABiBJsFKzLNl0I0x28
0W/CPja87eSnkeciUVQt//cfdJ/nZKUULqviZMh4DN+5XNgWY5PxkAq3v+0M4ovNJM2IQv6Age6U
6FFR//TgiEMyHj+oD32ZkpGf6sWpsWTtBpyqMGp7YULqHqTvQC/sbD6HnQtS+kEOLGMqrjpjQk+j
L/gH2tyxX6xuxJjzrD8j6qXGi1pQkhH37iA3UFlFWHixobyVPQFhbd/fsB1LLr+TSfsW4rO1H9ab
Fi/TkdbiG/DdbcCM5L7IYL4hbX8Cc0Xc/qseQaPKdIGcYYYJkz9OkuBMmU5thD0GrB5ljQj25wY6
aYEZpfBlyVKEa7qhFxJ+Owj2hcqFwl2dxOoS9KkmruSqe5eP/5IPWlTB9WvOqqehAdUX9g3W57iM
r3MxFVn7fckKGDHIJOKaIlp7PM+FRiC+jv+Uu4CzNFrcE3l3/hg7IHISUph9D/MtS3x8UvvNlGUV
M8fIIOmFZrit0Y0BicmBCECtT+gu6PEh68P9ki9mVxs73YzBjCqgtFtWZ/uxEZVcmpTzEUQ+HVZp
7ruX7ycTte/0EP/9AOKeXELJRLQpnHyi3/2PvbIJd1NO0ViH91dYRYOu2u4jV0Xk+3wqDxj2JdMf
kIcj7t3nm0OSbyPFNkj5PlRgPi8+tUVgrHlmOD+SYTrQI5Sr+g5e05EDubON0aPpdikWnHChSnrt
Crewkw7249xYhYuu8mUJvx+3mhd85YFZ/WlxtmkEDQFlaLeChkXSa19cdIIHXPDkFa6+IPYtNivf
+KizxJGbA57iH/uLUdhFeWreeQgmTYsePny22hahshwMbmtrTNwMxkKTcEBC22c/67Hpvq9NkEb6
tyFn0CgkYr3psMe3gSF6tpeDnyHBiZxu+oJW5VW4uj5zkFe+ljjl1jqS0tp5iQQ2JO62TbWXEUAp
j/Spc9Wmy9P0alyOlONofnlSvBvcgo6f/iImt6/+cf9QHNkwFGJFq0AxVV44K05Fn2M6iMVzaE02
ZZopzLlcsiiDoQ6vZPxzgrTGhqveKHD9bSzWCnJtYItOEc6fsJK7jADrqm9Cytpte2eq3ty91GeK
q0zQIv4PK1M4ME2ZDJ1Hf4SDvu9Vcfi9sreXKhd6+zSnGgRgJC8LTMj2wupngDda/8RgGI4ykg6+
Vm7FbKtJ1fGu5Ds+5u20wasxyCKkH5bZSiVRNDDECtAyo+XstXmw7DwFj173xfncHa+TET4b9wKB
/MJp/R7dNJjUJdEseJXIqWjHkx+SyU6EpWAbsaXV07YUP8AwxbEY/1oRQZBUwakqAx+lyu/wAOyj
x1tKVzouppj5KQGHfTubbJiCJFQGJ3REgriO5s/Lnfbuisllg7NlaZQrJvA1dEGAjYXK+ebRgSJq
8WFvfuYdTCPNbEPXL3A8lTQ22vP/6UhpPpe/PIgva5NOLvj4COTo3UAjnfSTRGwLbyYchakei3tm
f2X0UlOwvdD85ta/SF1s2jRHvdQ5j7K/00fG1dGBuHHCemWoYkLC4bGHRJQQEYiMvwJKVM3vOeCW
ET0JjxlxO9JbksvP3JnRSte9gytwWuHwihoiRDfflhPdPuXuREFPMY7UI2mc3TIlzQ6g0RViv9Ib
pnFB/vkU7TCEBBly+L4WYXdUXPUQIli++aT+fVtWpXYSZNBkEY+briRd95WFHMjjaWSzCyQulIRa
WXCgWgj6mqyQgqZN2dM2JMG6ERUIQdAEbdjcSvGfLkmtSjyYkKCsLtcf9KP6hKv+aSNN6zWlr+Vg
OkK/vfBIcsxSbaf8e2SEdF5QZ0ObgPimbMQgIrMBYvgQ/Ld9WZiDfijNR3X9chOHu0Rhs9N+Y53T
fE/jPOqKtSXYCx15ynLd04wLFgdIuQfzVflgyNvDugPO9dpdVb9Sb9h5+58eWlxtILssQcVwCni1
UFKO1fxLDHwXIK6r2GIVUejYmdrkbWlxqJZrPE0y+xjrf6Qvx2w9mlOZTs6LcDYqyP70XWuELbqz
byI5BpS+4XygBpRLE2vWfAmLypI5l/39knMpZzxKuzBN5A7iB/d7H4mzUpyXCaz6yaO5r02yKr2V
T6j5qZqft2vR/QNzmbs4gPye5pg8dnvIkZkQlKv24rD2dU2Kioz455MAwhAfrTi5D08r57PHrM+p
V9RcQ1OU7Ty00LftOZoWu833LvOWOjKvlVHZlLFDVY8iD+3TkMHMQ72ugAOKIwP5Bgo44Ryi/lnT
sRrHrWnfrT71PPB72ugsj1jlqfrKwbmGoUJFneaDIw2knLAkY/TfDXLumSBmu9kGmhqRRbpWc24I
9aYkU+IGvY7kLgb1qxYjMhVVMnO8h53xIr8T+jXYQGKBKXCVHQd0JM6vWeMRtlkRuj03AfBODs9N
4UMRLq9qbmucsahPpj9xcCTgczxQvKrQh2MBuwWQg9i8wTM2wGyarjB3LBFTFHIvcSNQB+5Xw3Qx
0BoI8f7xRUa1evZU+9WIJgBbfoVsu9BQ1nGYZhh7Ylzm+xCr2v8LJMHSlN35R6xdY2Huyfy1p9dh
8OcIdlMtmqKB5bWNk21PeUs2kqwCHnpktGBE0HNj1hJepASBXIbiS2qqjW+9BRO4OeYJADdp/WxJ
XT2e97tgPdLdF1VbDtl/JTzbtqXcKKBmL9oPe2yi0mm8tSgq/OOC6qb0I5bXaj8A+iBwCJhQPC2d
I3NUZAZ4NDpBcSVbb0bpFox6X9XFx3+L660TIO9wFk+zIjilj1Mjd/c5m6tQb0Sg8CbUoqzD1LZx
XVcCo0whSIKRLW7zVj6tpX3c3MJk1AaqLDYvPyy3UBjLwbn8fHuOpYVVzdL/D5naadzHft0Dzwll
Fu2EqVppksmrUkuzZ/MBE/s+u+yZM3jBpBb+V6NTzcJcYZWpPqv9+nhlqY3k1amfUL5lkTCDCB4U
IN4nyYhP2fszOURZZUyPrflxI9LvI2fQXTA0qB18ukffOUxYs9u2L27aApkmwSA4NgmWQSeLipGN
W9o6C696oWWSfFljifzazBNoDin/nUF85prJ70cY1DLcx4wQeLm1l179RnwHCqYOiAWPdOGxtwry
2xhGenWCkjS5FTuFKEHKlvBHVloLQzblLcn18Keqw1i/OpHjxlxgaBJCDcvKIM4WDSGma9Yp8twU
fdP3e/h/rnX5n/k5CRn2fqRGuPhvVXGINT8RHLOvwvZf7x2q00b9kY0OFwxTHL2sUcgOBmHKGWZi
jelfU+515/+Eat46BSow3C/tchiVCD+ytW7ohBoNOxDtOVaZlGVl4FmtetPBEkmSutNjEan5pcGU
RT1b2qSTUu5HBFUi61mFqpgnoHRGHWV2wfLV3+l6DwEBsH6634LUgbgDCkrXuzMKZQ4lvjpu4Wtb
IMsFKeRjqt+cu4XdDqb+BFWxsgGWuvDWI7s5uTXdcT+sunezDdMFegeU4jDllSkLmyTQBgIrctON
tcmSA2nScwLo+ECzmWh0v4UlGmZ9hN5XtQIxvVzmbbd6nuH9iwxEEkDCgjAXYhbl70n5yP8drKeY
58tbL4ZXQWgEQunpbGGV1QLRPEYNx/7rF4nIKLWktq8mHhR2f3KeVk2/v50KS4Vpw35W0djB0mIy
g0CRPIQ3hY8RGagaSVNKAIKBEo19P05aPtAOfHeBJc3opTJQrXGokq2K+NgG8SLmkOw7RYzQ+mwi
KfIMpERChsl0IgJxTBsysvJXPFCqyJ5so5X4nVC+jHFxmnL/ejSg1kr58vvNYUn43U9hHv7Vl+Rz
ItZvmPaP4bphs1x9J+7wuw8KAMHCR+aas1lgaCLq0HsWjGAD615DgMsgZ266XHU9sVsYUSNqfOzh
DtgnHrZpghjzFAg/pbvQZxOve4O1qXpPG2O7pbioc5L/BA3qtqEQocap9Htqa+iSJh8TE1UrTaqs
6JkC6SZXAUSViytRaUxVKMr0yY3kLpJ+zAfZyHoxsfgdmcKx7hdPIk/U7Dlp+9GsdAQ+etHhc+Zq
zGx9Cnx7/VBgoJmZLR9noWddxbOb/iJLOQOa1tOpVmUIPPifDAgQXkRDKKt0hdWhNKupysbXXyt8
GFVCARNu1OAGXm5Wmetr8afmYF74XZ4H25RlCEFwJuo9Gt76FFvgEqUPE2w6+rT+haXNdjC2LzqZ
mYCE496oKrRHK82eld209dHRrfybhhrVFYkdTHvsCldYuQnqyB7SXgiqEYJ18SrYVqIFqyNhhmE4
kGPgwlmkIOcuieGwvRM9uQryfuUNccyhbc186RW9vnJzfN73jRx8G3SFFT79kQY4F9WwsoxLWPfL
oL3Nv8dP5GcETWSd+MZk6GyukuWcAJfCcri6YpUH6rQaAVq1rsumwyIpS1+XePrPGRbDVOc5TbP6
+lFbqN38oKQuKDwyH+8JHSgHVrsoIr5HftDZQmObGw0mkyfWeHKM9jskpupBp1JZWNabH8z4wtpP
RNXxMtEIUh/+BJKModD3+96eyEoZAvY/ypUZYAeq39ozdOOzCjnQti3NWleKQnwSYnkLSjxsnjW9
Ou3yCG+eAVUUh85/pvYujOJJGgWxSFZR/CrxamsGSfhKr9PVVnm+3nT9xWN85L1LpUdQ9Ov/W9at
8a9szpOPLNc0YXcI6Nz/807yVjmoyF2sA6bSywaOBpjLuLH3CIhLBY4ZuTYvPRJcSJQq5w11toXq
lwgt7xtxN+d4qrgq+pAURbP3lgzfuDVBeiZkfzG2E8JX6T6YnUenamwipQjl9Pe/yMqs+stE9NxZ
k1VBZkzhYuwc40wFICeCXAdPJqpWCluEJyt7m4wq+xCfZSLLtzxIj2dC27YuuUYp7jVKts5tOBEx
WdSIUZ7PZEpucS6x8unUVxi1rudBbrKSD/ZHRj7CJvLvmcH9oypO38sVRYQyDnWIq2AP+bYyL64b
0iFr0B+VfOKSYgEP6EVLsycOLfnzKQhGXDH5OFSdJ8V4KOlJdcJsbTee2u8Pz1gFYWjIQioRVlll
VbKpIeCrxo/IV5dTrAnCt7tciCS1K1U9yEQ2M2LFUVsyx6LvEBP2MnPLqDwHrpjZtJv8lIYfsJuC
sX5x8GJD9Xx4F0PT7XnGNKlvuIpP5vNmKg6mKdzCc+QRWwM3/1pHjTIFefH7+pfSSOBK0KDl4EiO
BB6bO9xQXFOes1nOqrK9PNOL6bBi0y+M6rl7MPgr0J9roYj11vF1otb1fcFDCUZpnWkZ0Q3h8hS6
l93EFYq96dqT9PVuZrrNg9OC31oQCdFruLfq3qAOqKDSV6U2iaN4VtCk3ya+DMcUvMezh02tGXGW
mmGdX+jIWuKGk+x7HpG8GSWnzMypR1Fw3C9KPexXNGkMb4RD0UfPH3nf8l+MHdT9muqjLj2/pyRF
YD79Q0ROPbV0NXKtJhmyVzVWc65sMBJRO7DGwr65EHhD6ppBx2wlZa4JZvysbKyExOfk75M4Iy0t
GLj2luxTwscGi4a0IRzSGdFhOlzchzogDVL/xWkR25B6lljWGlxI3xNHS3zodaiSXRtnEU+O8O6o
RkemrrFvFkuFrntv7ZDDZc8iZVBAtEVVK2gyngVQZQ7nSG1X5hRnVl9aYfMzKfUCZqOMHtCzEj8g
07xRqEGaM6PM0MWys7WCIWYvxQzEz9AjX+E/OQiITHfkaiuOtjKvyzs5ixlVm8rGYo1jFczdEuXG
d7X+sblBR8PbjRQd2VALdoQ7mIwpScEYkhckhzigqZx1kHOf+5fVPMg8T6cGHX4Q5Hq7Z6+iuoLw
z/oV6xxr1vQvowAcbAghmJejhChvMnq4jvePl8HsX5IJ2htBu5CM4WAyvZndc3/JJfzUsH4Tsa2O
9QFbphufMCr8CfDSPj/SZiNSj3MWjNrBoDVNgvXtKbwAf2lJ5kCOcwQ9o1FRtub3GUulkean1/Af
eMrCNwq2wBz9NFwpeZT03PePfL0xqWaiVBEFwmPzHHoOOFMSSlIW2l70im1sOLz6MgyHt9JT8QB1
dWIzthmOWfj+FuCVztW3hJK2YJAM+AT2n+eA68VgJNkVC29xv+0aDgBJEUNVZV/sMS0b/9WBJ/vH
3UoidKbXS2z0lgfNdV+1/C9vFlvP2l0vnqn9En/g73vI02Dl2cyWNVOXDHAPEUHDcmqpUV55XDjp
yvAyQlROhVY/r+jiYiSbPCai1nYfcCIfMHcGWb/3hlwabg8sbLcYAuIhh18/6hvdEdGCnvgRfo36
ZyYxB61u/VHpVS+QbGu1NB345PUD4MRZ7AnIpJ1Jfbo9b6gay73sF8ByFuW6cmfQvIk+xR2pywnH
CTiZEl2BwrDsBkSzO9L6TJD87YBwa4TtkhTWUBKMKp5NT4kTLg1pvdneQRqCYViyyZNdeW4TRQel
8h0CdMln/+XjZCmaMDh/6ib+SPGNxVs2SJpHce6Rl3BsjECLhLDUJ/NTJXT4AB9JzVqbQ04jmbei
41Y9JljiY0sQBNlmnVgwX+DXT7D58/HphoOUbEWfLPHSsS5xSscAvV6IY8OlgKjfg8wCrNe2XGU0
21LuOa2/OLCIk4EGQSlhCQWkzPEg07juZCGp053QrteSv7wO/s0xFQZwX8sJZOxkIlRK6Tjx2TGx
9oWXl3CTT+L6lp1numtyjB48mhQ4A/glcXDE/xKRiuqz3HXoj5kdIo4l4s3L+dyiab59+GIqEUMO
cdp1iPfKwhpaREMjddpddcglQ4GRvfPLwCGcC2tR9Psq+bamgJmPOBPKtzbm2caLVoWNIE65F7Wo
3sti5oVwl+tQSpwL6AfZ/1UoZTrmVsbaq45DAQPWEaHGSsJapcV6ldahLiGcwCh6HDlSjo2hmbAn
+a0LQ5vQXcSGHxFVlBZqDPEF/GtvpNus+MQh7wUi8SzxWznMJO8/a9wauCmdjZRyYvG8JpW3SYs7
81eIDhw4fB9ngzJVZM9gVfPozArP45ihWvz717r5e0BxYlWIrbCWTPT3Fkxk3K+6EKJ73aSUpLuX
zdR23xDDIwxOtKq0deM9wlA43nh+Frt4hAY48npPdyoTlCqOb+f04FWwJzHzSyp06tzh2vC6IZhy
B0bn1JiWHVf6SzRWd4DEAMERlYp935WM2kVQyWQql25UHcZGL8H5ITlaEAtwK9tB7TLVRoSzYc7b
RLvPdB4uB2hwOLgzr4xoEq4FWiM46GdZf0mf29g52FqlHY7jVvvFD2MUVE6ADkC3pp+kxaxvHcRF
me2srZLwoMIRzvX1Af6qxsf4PCrUL+H00S1nqtbSfvYVE8HlpSElLqhWs2zGYTHC8Cw0yjF7LXFM
yH/G866PUvp9Ee8zDcjMVWC8Cmxiih7G/rczuZz0dWArm46ZhKffgD/KGZI4RsceyHekXEwTvtQH
qX5ZHDMOIdpgRLE2SErG62Kb3chjoioBMs+iCi04hirlVGq4BT7Fb/Sy231CnxX4tA0P5coa3yCm
xaPchPK2oNdpHNz1XtdO939OHi7mvZMbT3yty7UCI1qWDzbTr2TwcKYYEVVuHeXxDoq7D431/EwF
KL3h6Ev1pxsDg0frpwqQotU9OKOU9PRXOm6VlaoxZEDIakkW0ZATnk9hWEjqT9lpO3WXmBpc2jOA
mnnY9e3muCQU4MII/uYQQ1Do6wt9Gk1E5b5VUsUTW9S3dFYvZ42W1hP58uAf+OWyfs4buvjI5nOj
7JeT4v3dqDQaxH+bLRPq/R74pSFr/YlzlKRG+JiEbWzA6f5VzQtsEHPZYCDtZBvQTgC2ijAY7nZL
WSJWLzF30utozid4smRyKVm6drkUYdGeI6EZf322vb6w77Dm1iQwxWcZOT0OFcn2PhrtZRPUUqHG
0nGFRRZjvqJ661k+SIjMB71xdhj0INPBjygVduTClUNTzlX52zrVMk4o+kblr/0gzJNP7EIT6wj3
O9OtMfkloRIaS3+2dSygI7xYiuOuG6B/jz6CFk9EFlFiEDn/XgQnnvEvuEDmU7mjjK1xLkxSIWMi
9jC0NWM6d1knfoJeq2FPij9FtuNiptBvHfnPJjtDVZqO57bEKrDZgcxDZ2ulQf2HLxBQrsEBf3aZ
VqNv3RCgQtyO9tyhZ/IfZcc7fBBvAiWpyiZnAIAQyDqmwYVy7+YkijRS4ZZGy/N4G/Y2s+HrxD5z
545iTWAiIIhB3eraTd+1IPsrXxeNkHfyNMK9t86dAdjUjtZd/X6cqP1hXX5t8VrdoUv88Z+Tx9d5
SloCrj8L+MBLajM6j1MkmpEXk4r2jtexn8eru7QsgvbqtTkDo4ZdctjtWrd4alHC14ENxGSNTB7G
RnAUwd9DXLbqR07sQh/6s96fFzjx4ensjJhlLnrrsKwtkVW7gg9G56JThfmQlmdhfoRU8qorp3S2
sOmJVEsaW1l+ShYNAEiDjF0C7NZnWiP9l8+MPRvE1cipltkFR9XgbUw+vPAhUMJZlPYs+isTj+mI
4oxgnhqm09PjNMPiw7Ni874sjBdPbhhuuVil4h4rTCkge90p9fS75raZTFq6L3xcGNgOpJNfnqww
P8vhsJ0QvAa+f6qfHYnuRE0vFaebA7Qux/8LblfQS2PmDrAXIDt6m7739cdsm0cuF4j4ZT9rIn3C
BlCwsmcKlLHV4FRYYhoVo9bOkdWiR/y+JGiZ1oYjF4BOBKqPIYaspDH2N2tqNaVeSZ1KwnK76deN
V3DJJdBa54HTjJZQ9LJfaEeXK3xUSgHmo1PTb+ofKjcu/4jluokjliX4xgXowB7HM4apN/47dX9Z
wzZGnhJqVHNlVVBZvq0WxstcG+waeypOx9AoIA5ubScYGRwkdpTdzVTT0HhqrraSKop/gkm5tPno
jps4F25MU8a/Wq94o4e1xW14i8+7z7FdriBkBDfPE7zSyF7rcqfhR67Wsp+y5z7XYuytgJG3PxvN
D3myWhXHZ5CUonta2P1s89MGeN+2yAyrZSJlnbOZvsSOrl5AcEUumMN6X0luoAo8Jjtfs/xJEMwQ
/Zz5yq8cUcZTo/K8q5IQuaUdGuRFvHHYKNZZgFmfISmAJeZfuQfxYhr7BIictOgkXCrcI+N7Urrk
10pp/13ISipBowBhkAwo2YgzcN+t7/IJ/zh6OZGG18MOdCiVPj+KN5NlIuRbl/Zn5RPo7ILef4a3
dedZgOpTrttjyRDXptR9RVIbM/VXGyYcNYyaBGacDzbrleXq5CzlodkhL/aJe9MoCx3JI6iIjtjn
E8OA48R/Qp60EDoju5vfAlySAv/zlfMay2lz8nfv4KveI3V/gg4aWodwxqU5FiLNmkIhiJggh1sI
4h8lN9SZfMBIZrU7u4jLnV2CvM0stwYqaOsqFfQks5NNQcZfvU5AjLD6rAETdJvn3CQ6qNmdK+Ie
9OzLHfqF2eG9HDkQU+Iknd2RRq+Fet7jyWLS2SJlna8uniuLFGOjPqv4+7QNqyqqF5oTw6swIYKf
meOQhnVLtWovZ3EIr8Woue5GZn9GKQGZCSmFzJ8sX3JtIgqCOeHaiG/nVNlivO8lRXVPNUd4xIEZ
PtGP9VC9jhj3S4EZUf8V2Q+4XqjtpiNqHftUrToIOUCQEqgrvt3NQ+nk4TIKLYkAFHR+ikSyF/ba
m0pJ52hZabVUXJUe8udsZSjx16N69YNLAirWdzPrVVc+/1PRdfOn9D4JJdOy/w0ZBqlGZ+Dtv6QC
A+vg92Ty94iRC2S3eD1Tm3PBad4j64V0Pr1KNCCfYzdNpovfZKUdYt6tZdLefxMVHe3kSbqSs3rF
rnjK517zhYskCc+/Afe1mMk07fIi+sfPbOPSpj8G595baVkQEtrgdMM9kwjQyCoGe8sVgGjDJH2l
yw6KOw5Xtm6bNqRZmmWa2T9DKSvWLJw65rplScj+2skFjoy3a2euMp1uZFVQ+78U3I27mpmsEwuT
84tjN4hlJPO93I9FHDlsqf6s3IxmXMAe6Rxv6+aCHMsHkxUdyCQgzCXiHmSEYkaUVSYN/t8pJyY7
064EqGddgPqHrhivah/34ttZygLm7YHkq7XGkKaqHXTTPiFZ/+dtW1XzcuRFlSy8USYxwrhymwca
y/cs+Q1g6sqny3S57dDKiMIKMcuD36/dKp2aZzVekUtFGnjg2R1YbPu7ugNbCYAKL8C8n3KQj1/6
pmnFTyxqrHGyZohPDxpmM7m5f+1rDs8Cp1ZvAZRkg9h44VMS+Eabc7MqaGcpVMaFiI6KjjPa0m80
BjakeqMyAu2LrzKqLA8hpqkbB1YNQo2N1bunE/zEVx6hZZJI6eUlP1CAcBdzfQqCM1wQStL3lwRc
SexIit0gcGG3KWq434p4TX7DkjGPfszFEJ5aoB8iX0NvwC3OrI+7WeEq072sossuO3d9d0FBPONs
QwLfi00vH3rSkD79F0/YO1FHZquC/hFyUUcb4tbSJoRad75NsfgayncIcDbru7C/ActSmSUlacij
G9pLQQVPdWNyciDxUPIfsNcTlbSaQb5of1Ju+8XmqHM2RQhUpYrVEQlt5ixtZZj8Tgko4Ru9LxJq
nrBBeuOBJGfaDC6M647/YlJyn4YiNw5wx67AA2PwGNZFNummTaVhpu2bbd27aQouM5AqFxni9ZLo
FlvOcMH0LP9oIwC7xc2+7uC/0D5CZPcuF1OEHJwcQJ9lG5q6yD7TEQ93vVtmvIN8Jm4FpsbEE0fQ
MZbUDvW+4z7qg5Iqjlgfs3vsthmML1acvgdCbpLTZ8AL1ShXcbo3TJjrfej4K/oYK+zyfwg4WYs0
sUdZRpTFyvFkadfiWtxslTHwFRcVdODNgfHF8xNNEgwHNMWG4gPFpN2CzlwwkiO7z9MccI66eXB7
JNNCoJNSa/wgfGkoXg0Q9EyLICspMDDVUxMnS7emCcvTq7wpUBtmWYSwbfa/A1rUl0AR7PxD2RPH
VpNWzpG0yLZJEd8UIpCs2lkJSF9gDjQhSLX9BKC2KwrwH0KT9rKV23fVVfXxfIMVu5nCg9l2Hu+p
wkD/GCEFDb3WZ+xYCY5ktCMZxuWTdpxK/YEGDjOIzoUeUqLscFEILfMtkKses4yQDDRx1GtYwvjr
6DuIDBwUgBK0zswxahWs6/wulLF/m8KU2/cj4y90Jl/iiFT737opby8HZ5eA08yVS79aeXhCVDno
hXqjB0Jq8Krj4aHF1DiHOi+f2VbudXR1XesxEyKwY3Gap10ad6i8tUpWPTg+YI7GFCLn7q48CLx0
HPI5QLwq/5ZGwxpmGfNjO806wGNh0EHwoW75mq0o9xndz+TX4vBVSD/qdHb95Rh2nIMl8b+oOhoU
QTVRljMbEsjkj506+tKxXD268aGB4LyyGbOVKnT+525u2WHd8QfMa7io/WzKy6+BkXgss/QGvS3M
20mjBM/JQxLtESqxNhQfiU1Ln/oNTCcDDfpz7/+So4C0DOYzSMSItUGQS4FfLurTj0NXI2d1Yzut
MNi7yQnqP2nEpnGKHZMxgnL3mp7KVoAbtEnszhHMiGumwHZyVY3toXDCtwB/AL1/Ye9d1uoHygRi
QaR/NAWnE9Ta8peMnevlnB1XYf1J2UM1mxlytCw3vy3xl2bCJKXSPBLgLrT7G5RhwYfBPMnW+jKT
QY7Gbcp+BH58v8O6xxAAXwIG2SRyxui7TglaUkB0Z48mSgZjTJgeI9KUHyCubySqDRJth/YhGQCk
E1vYBxSBiRvSa1u3g6OfqkEV7SyiHMK3TdgeTJ1rhZaJ3KlWLRyJydoWpR5db6CIF87Kk6Dgeu4v
qL0CtmchzZ91Qtu8IGjUhjLpuJ/2n5OTCWUEU4XFdtF8uMNN2+wyhgFa+6ZrL7LJr8lZ6g2uQqVA
CV2qmwQ0QKzwa5whbZ2+u+pIcqeuDOybYZiHY9xqhntF0TNaVsyiihghTludzJRMf4lrh8uzPOL5
2PAgK0w5kojqIccpdZH133T81KpAdyBT7tJ2w5XoYwklodr91IVhYQ2rtYiDK/PY1lWiEgl2OPyn
3xw7d/OF4RVxIieeGvnIAHDqEB9W3or+zRrBm5jaWgPySV/oM5B6FX8EsEjlcRY+hFXVuniY/pUc
nbvdX+vt0fxKOae/PsQrd26ttv6tu+mpBkjaTCu/ZGVVRGV/lzmIihzIyzJJXZIwrZx78KoYDPuZ
JJ2EgDoxsXRq/s8Hgk+V2EzaHi1wcE2u2VzZcdezjrvyqnko0xwCS/cK/5AhnOluXc0prhpt1TP/
Rn71yQqmVlO7KyUrtJsQsJcnTrImFAtjpxTXoDDA2ZW4Ni9Vh29JYP8I9fP/ZufNk+UBAHi3Kjma
Ogysz7kAVTRkRrh/1jXOFI4cAXivD47fLgeRJEyTVWnJH+SYwwXfVFIooGzNfkK7AQalUEOxInrk
uVpXtH3u6Y1xvOt/VaECe8ajjx8P2EPrDZskTM9N5xUSsX8rdEEbRHe1IZo838IZ3ThpD3uAiHn9
hYNl8kTieztl1oyj5eXCIkucCEosgT7NNpnGFb84dzg+fHi6hVtjwjiIIuPM9Vkcv9Y9lyIeAAMH
FY5X1J+lETlxAAYiHqDxRNFNXT4+FthGTJjKJImWFxPdrefFGZkVRigasJOgbvVXzAtMkOYHhGbX
PEqyPcpfnKSWavNp6epHnv2CjDJQLxUZ0UzZX9OnfJQRQP4Z54dTHUHKgPcM3/St6At7u1XEnu5K
eB72y1xDXOkuYNaDB+E8BJQtoTjpLB+pJjKA80RYNF83IGX6U+7VoTTkq3gEcnaqfQZKo16pP4Xr
pgmSeqnRs9no+hMmiL/KK1hBMCdOEiK51PCDtstDcyrcT6ADmXBiPY3gVgPZvqjw5WAt+u/0XZaC
oMqNo0xGUhg8/kKshta4HasPQHkI1K7fK/N3PHeIFqs8BQoLYTLfo4KV/5sHN2edygn1evBTN1Dl
os8Rz3bGWM2G2I+bs7LLSF9jpXCiAeWlBKMUPotY2Ebtcpmvx4QqUZzY1BtykKAlpwZF+jcnq8cN
G1L/xtPnURHqUq4kfFPyHfn9vaEcATCtIi5IZVR+e8FOIX16vdFg+AWbIEVB+OSiZLU+dSXqV8a/
xCknJgKjkQyu9mGsSNvCWkU5JsFoT/4NdRi0PrUdo8hy7Jl1XFgsqRevue3Dbt/hirbauuQXNuZw
sEie4YOjDn1JmXcfqf1PzSj2xlLQwWuswv1UoXJ0wWecLBidM3lsGA5mBcK01SRTILCPANPa0SxD
0q4dLBBcnK10osVXPM1vIm4QSRXXYCjl7FU8VE0x5otzkLyP71bnS/JJg2qEsbmUnRgXSUNRDGRU
IDmpMA06kQI4xsYl6TNkAZj7AWRo88aNpRqZtQG7wj6qki40zpma90j+iPU+c0W/HKUE53Cqn/Zb
FqZ9gWyGfs8m+vAKvXwQ9peholJuqqJ9b5gfVYmH00t+Vk21uP+YFDiK6kP0Rxuhw1CqATpUpoZp
OT56qLgqiEnQFssAz/Xvo8sxzlUR/yEOnlvBQDaRHJF9Q2Jrb5o0XeLHeknKq1nLJ3WIn8xrU2hS
qZL49Ic9l5y0KD/aKbEoI+kdnoKpByGsK/wz2My0PhxebYnUaNEDJjn1Spb8dQhYIwt6GFBmMOog
s1Ulet6Ee1mslEX6HXvRaMdgwPa+Py6qAdJUXXaKVsm3S6ma4p6Lg5j1tXwoF5w5ankDYHmZeznz
sxDjATBVCnYr7yumfUvFAbR1wMiVLeGhIEGx8y0wa6L3FWE8k9ssOvrSIgle8oULlVI/C5zgt9XL
yz+tXHwXhfTyrQflmwIAAon/3OAupI7X50huyDdjOpfFrpDfjU8gvH1fsQ5xnNeq1PZbekkj22A4
K0B7/6x5BbzAtzIIm8qLswe+hmQP1kMfF2xFLCmVEBjUDCQW8wWXRbnLu9K+VtNQfDzU0RwimyQA
3p4DH6EnPen5uKcaeWvTQnlobYCQUlasm1b+RJtHZilD3g8Df3eyRBXmgIiJ2On08TlGQ6ST/S71
2b2A4cJqqke1N//847XWwKqm10k9HjKXBmGIk4rLo2s0X7ldTt6o+48Vqk0PhXPmXv9wtamLXvRj
PgZ8v5Gk+BmbHmSujDmHNcnnkr1GPx//qh80YeMFtf8XqVmJM80KXu1LJC2VxcJ7Bg6UR0YeNvR0
bPELPZb46g1wFi+r7RgzlJDM7ZJnPucwZO/ZhgwHaCQBrwtfqd2cFoAaykN3ZLkSaLWf9vqpeLod
/DKVtt/zJDT0czaCbEo3xIAbzUq+airtsEi32eeSv8rAyrdvFJORocPMgvcvL0e3HKV+Pq+ROOIq
hpmbKM97VCQ0QHomwrCqCubT9U6Ot4jJP7KuJfGPAZxRzxjLTmo7M2eVYFG5Bt39QS+bl8T+zpJu
jN2wGDiz6rxsAA/Wzh9wvjU7mrZ+dw/iMgjq/rKg8b/bQqt3r3ZOK23UCrlUjl8PyyllMZK/Huy4
I2PuuyXOiAl/fAKrg3KS55Wf0Elp2eAuZJkjeiEw7AJs12gMUN5PbavNxWdq3zfPQo9V72IrUmqD
wxFCOwkQfB4F+APTkXd5ZZiHR/Hsm3fAR/N1Q1HEh8hOEMS+B/gDTBXbf5a5kl7LoY3/4haSfaZp
W4n6BFPk1/9FQoDqYX/OwItQzGyQC8Zma2ZAC3/7aMYSVTqYOMOdxIvcKxgNO3YVFxvJU1PRphVG
8FMYTBZ1qLXlo843Ou9Lw1+0pYQ1hilsbgh32d8/J8rXG9+A0d+gf2pfvkJPY+1+xelvL2KanUpb
ukbTe0New0Wvknr9FjHXJp/2r0EV30edG1Rg03NgFuQljuFMW9wjK2zC+3ozKzEjM7Ivi9LFSryY
kqd1gYgbUKqrjSMQNHEOFlrYn8awLld9L5qWr4fXTU1v5IOPk1yBFF62FGN2MZyQprfrZ4hmlEQM
7TJPd4bPu4bF6ohUxD3xvYKTjovVQOINDvADRATs8Dtr0VuxT2SAP6pWh2Z57zR0/4Yk8Lhl3e1e
vAZxygo0PMhBh7Wsc1urWbbFblrQWI/DWS0/DqwmAmTZGBYjJTP6ELlqc/vKTx17aA/iCbjJJB+R
K8reoMm206/hWnQDtcdjbCBLybrcXyOcaRw99e+8+f58JmVg2fWqUkoTK+rkv+UrSTx0Ovt7DtbK
JbLAyN5GY7mYlkWfR/Kkb6OpcEiO5NS7vzI0YDkyp1MG/faHtzzyHM2PmLiC/HkajguXwUvPRug+
OiklViNCiFYnHB7glgvNfCAdZ++25U3rOtJV6KZQkTwAgV+NIrbMebG+xyCu+1ikKOCqgUUvfQN0
FKCq5mY7UYAQ2BSXLwnhwLFe3/5gL2BQBTBSEb15C3n7SWWrzl0dBUQ4eUV2zu+WKCR8ImkC+/cE
DpRevNxqcem6soVgNbcqOqiWFiv0DUQAoThgvWx6WjOXlTnQvXGEOUTQRscp39NgNJV+/pnVUlrk
fRWuN/yIRABgOZf/ot/wTJOdcC8rAg+6fcDjUubc0KaMZm24+dyRgfbwrEJOyN97ots0yC3P7Od4
FjBDM/DBqccdWsvOnQN55eyzASjK8aEZpEcphp/tV9xs2I6s4JL7kvQKglCoBase4813Bx2ZegGI
wGWjAia+rQ6YKW8HXADb8PzFWNAyFsfb1b675UCJaRwk8fgtDvdwPTRJfbOzKuZ6O0C+hJrbcFPV
sVIhmMH3jmOt4F+uzLq3SJMNs47jNp1NyR52GoAPollTBwT/jVLA0CNEytQwPH7CCbfX9ftWXsYI
1HWtfnyn/BI49DuPT+0pElysixdklrLcKS/RPAHmazBgtJKAdjF1rxghE2pGJ/rM7lt0J6K6xyaU
TO/HD560fmGr3TgkK8mNrhYO/+iHM+9QguYqCk1jWJT4hVjAWZes+aIzW+c+ZDDion178NRzU3Lj
GQVx6uufBnHpdsKTrgQdoXJnWNb8M/BIqw/MfZc1nyOe9EA9Aho5oPpSzCXLwqreHDPwS+HVgnaT
SAiTLu/qxG3CMwKTE0y1AWAIiMBPatrUIMWJAurnYc2r74Rp5d8dITigMmHQ3k4kSF6ysa9Kvswx
Z/VKCihxoDs7oqZ52hYSQ3UQjBdf7EuvdDVblMhpEKu8+5forNCHyk3wNpTSTZabSyfKuXsvxaBM
iU46YTzchiiJnLisylCKkPcACs7tvAJ6cXacZgVFtsFqM8f3b2oz4VqqqMvtq9X+akwD39QAGXmj
ZbnoMd2DN4yjvR9ghPwb8u6sAKfm2JAbnMvfCDJ+DsXjKDF7mqKNmhqKYcJBmzq1cncxresWh6v5
XIEqAcHcg5XcRXD5ygTBbUJpBat8eOqLIqXHtvZeGi6kuFzN/jDEZmxjxOXMLrkg1gQjO9YVaTuR
zrVieOEqzbJVcfJ6n78sA7Fs5C7G5B6QE/ueNPx/NXF0uPVpV2KPoPFihJtntCKENFBckVR+VKOc
91WMiFBtgTZxQVjGYB1UlS0ZzahDk/eYqfOwOS2oGKQIaoVeIGW04QqrF5WSrt55KEVm6vcnBaWb
78BP/+EetMIRi3y+aUk1hZuS+FUrugJXOr8tkSkAprric5U7FnIhgngkrm2GuK6BgXXbmBBssU1N
V25gCl4j2Z8VAh56iwf7ZKuXMVEHdqi8T+juqzjZ1WirMnSadKxUugPRDL51J/foIeOOuzBMVQuO
SqcmnpIiHtjE/gITYvIJRq5ZsOQt8jPQzeIL79jWcMFDsY5x9GZ3h9b8pwbXWAa7s2RMb9rjm4P5
BfbXvZCzpeeGrY73Xf2dg2oi+dFZDo3zb3kexVqRxOasMgOoNWdN17X4yCt4WHeNS0AkOwte0zqm
FzaKIXgbgah3VRZ06FrksZDdwkSMlW0SeDiypqY6Zp51mJQvpVqeHRaCfHZmMPbKSlMhXWAKg6sG
GQfAmDT6rEZTjxGfGw7v3oHP/0hiPxMSJmsNz2VlkJ914DTQA7SAOtutIuCX+e27iu2ZFeCz9JBo
WVOA0JA14J+zUV6ykgLaGgfxJchPvUPM5dMufMrzkusJkLyo97GvssF9adLq67Y25jPFXsotnKSr
39PZERjsuII6w8oYVqcrs4L3Pr3wU+ZFpmEhPLAJf+1rKhdUoq0hKWOAUX/vgpEeyuOOwjmNB98M
WIaDRxkjByb4qwwVy7CMcrIcsk21LDKhMjTLfjtmPDbktgxqDDKPKf4CqFKYptlNkQcjjbThkVAk
ADPdyr92cgfrVkIcdzXxjmibwk/osC595WDjH5uZR294CSV2aCazgKnh4dq32Wcq24yNICgax6OU
eqQdUZ8BlyRtoV+taq5RyBz2GFNkG6N+jcBSS1IXsgi6ZekhfCxhWd3FfXKVP0X9ojssGxPv7bsw
B0KQycZHk/CDa+87zKoOON7z7XzJ0wDI5VEdvkc+oGK6SRjMtdhdsI8CvmuLAJn1mesn15dcC/Kq
kWoH1Nmh+XWaiTg5khkNEUQaG8mtyAVoicxzC7FLBkcHGk50U9Us9HHJ0bVVYDr0AcB1cKDsUMZh
X5cPNnZ/kRFMDp0DJss9CoFPHTP/iu0fHnVLH0OY1UoMBceTfZj4g1nAmot49r5djYZR3U/FvC1e
H+3mQxQ70TfGdnOe/HVIWrUk9Fq6TcCf0IwC7lxnwSmgQJE5qT6L3FupK1XjAqqk+lmixVvEgtUw
AgMW6Ep66TcrBXWSSUZACwC49N9hhDZM4nkQzw+mRXGncqmcPasTUBJdahwCFVXxJmV40UiNiHTH
QFSmngEf5aNRW4PFahG+oONNCFKClBxmq8BgUAJZTPL5Z1YiletYr3pKKwaO/n6IpYNqqwcYft9a
tTo9gJYTmnCkMh6ZuaxPfgWx5F/yz/ZR4AYy7amVmtvjcN4K097+XgUxD4MGMeWCTbqIiGqok1G+
Lp7ahq9hHTwUbIh2/gJiGto/5krRt2tyT7VQuvv0M26qGb3oqreW5M8kGVLlfRFFhbdtSqwtXqdx
zHfCE55E2bWYE6JUna+EfgSykdd3EtxcFkXMZH5rCbW2mj+I6a52hYcnKZUT6qbeaU2QHH7C8uBm
doMk749gaY57RHh26x/0TgPCwhKTUcFEaAQgTZ72mY2PKh0NzphteMb5Za/r4/fwgnzfV199s2tt
XIfkrrmB25jrNEdJNJ0MNTeT0PKvvavwJzN8tg0DpudNWfUtInxBVYmQ/hXQ7XMVaFYF8b8mvcJh
UC2ez9oS0bs1lW5SD5JJwILmgVpvcC5a99ajO1pY1edRa0nXhwggQ9oaNzIVNiIJbPPzz9GbUJjS
NNVx/WZIGFcMiAtqg0Ch6pUsSvPTpWeIu9Gmdeiqeja/16FJtOsSYZgLmB47ZsQsQYwT14blFa6w
7+VIjOEcHTjT7CL5frrnZhG0hAEfXK03GCpBQv4Z3zYL2YobDwuWzaTqTitF02gE+DNz/qxEHhLd
UCMFET633PwwF8MGsE/xbKBimieKi9zHe1zNgr3M2rv611v9P2FFCvxpV2A4UcOSFU7Bx1jw8wLV
4iIaeheSvtm6Ohgxch0Fl2pkzDYsFlgDW76juHUQFT+1vcR7CJD8MgYS0hgsM9U/X0nArpKfQMMY
m2oqiwe7i7Xul0QvPuPkoHsEH7pONSiSQzmUiCxyaNEItFcztjfYOLlbGHjmdJMtwmCjaWXB6w95
wmLdwLP7iG7NSnLnwd0ZCoD4C7wchFKi5XCBTFJBkGhBNjqbKGpp8Ams6R0kQm1/YXIpFEw3rSVM
DZfbzjNTDHFAIOCnKOnk4pHyBz6gZ55SGumcFYvSV12qkcgdHtRW/YfT8EGNX5whvAfgxKnTn+1L
FIFaRJrxPjuyGNJ30P4p2nYeMx96v8WtwfnnJwCTtb/xckYA8/Pt6oR1eaZdXYj8ItY6hivEOhQN
Zx3FI22Y1ipsh2msHBSO4XfkZCQ9+2IUscPifAoCk9F921zOyYBkSPMpYZqrISXXJYgRlEN4xttb
9V++cDUSRzZvicfsjq+FHQ0NlHhU6JIo7zH80IfQjS68RB+1STcaGYouaR6sklpkxHya1HfGmjSV
ZloDticcDUO/nUHhP1pVK0YE5mPyctiHKORUPKmEmtsx8uKcM0LvJ8mFR0lBdMRShuf2WPPUr3Zc
6dHlLJya+HzWKpi4Kt3bkMdECbOJxhpQEyPC7hBtAp0ehEsdFTi7Yy3XPRb/0p6VYLucn6B8rVOr
LMW4Lq1Ty/O9dkhaQKwi8tIl+zvG74IL1pysgvZ5TdFM/xqEhWDqufbK+7w9jtF81r+IqyBLQpKz
47YplR20hrPh0OFxCiHmJKbt94NDUUBC9GdadwYwtqmsb6d3q1aubCX6kcNBztcsbMAckyfIRPcQ
RP4Nr4hhj0vKXpI7YLNvpGM1G4QVatMspMoeYS/ywpCY/LwXui3eK6U0LXr9XfpZQODqoRPg/8ly
biKAItVgme+eZklB0arRkxjge0lx7byfmzL/iY1qlbyDtNh/fR63ps9l+yH0G4agTtKRyjFnvc0L
U2jZRn/3NdFShWSddEk8u+bcGojSOyrc7gKquHG6M+2A0AWmv3Eun2+wC85eBxTB5Fnk6lFHN86s
9GY1oZZjx6CptuV1ESk/b8zIJVbZ0LnQ9jwsDR+qBWlSjBdX8ls6NubZlOqahkeIgNOfhXSbqeIM
C772Bdyfx0BHk8D92mpCdt6OsJq5xKH+j6iHDVNC2oPVov9P8hSJg+ZC+5JD6UHUd6dsJE1fSV/K
FaJ5rb/In+Omwu75d/i+XvL0CHyuGqydHfmBxsSp/W5UlGrpRG/gjfDkBKHlBQkDgQdvYANxTp/N
ilpXJDiiIiwCl8E/cc66m4EmG9UJZBD+3ukRzEVK7bMomAcMr20vSUw/PjQT+sbvQz8LLx7eHhSN
4AQJ6xgxALhcfCOrtIpC6ZTbsEe1jMov6gEjOzdqT2r8jpy714mQcd0Bnk4u2rolQ+dRedeWvCZk
5qNbUvQs9IO3ugg+iGR6Bqm+wuBqsBX4XgXbSC10SjbbWu2OmOkJj+pWtK15knnGLWFyCcW+UBM8
81qM8CgPqdaF3Q7cv298li/u0Xqdv0y1zDG1RpSTP/c8veOf6GBJR6SoUGsv8D4e0M9a/z5/au9w
r6xV6etFYojGDjFJWaMwG0qXbvHGAzggp86KP5W9piyBwRs/fxqykDH1ZE4eR30mrXgAdt3kzrji
90cs9e+/y6nq5/oNISpfxmFf1EFGW4HsZIxnvuivUaa2jHijYEnCPro4Wzr9J6x1h3RtTrH3STJ+
8DZlih0oaeCjXeOgQsW+pAX6rAlQu+K3tcAaYolNx9fA/y3wkrW14UFLs9l2QuC51ESgPK7uP4f+
B7AtNRd7t7nw1Pijuf4lnppzmbe045u2WG1v4e/HdHopPTf7/oXyPMh8mG4QaFNLEzdaAwWrhpkL
pT/M88+9ljLfbhupcIzGbaco9FsaU8se28pfoWHWlJBZMi4GfwMkZsUdjmFk9pauNbC+7uzAVQhY
F7Sb1D+hDk/tzHYd3odQRNrHdQ7Gm78Q/eOw4rMiYqBk71Xjv6ykkAubG+gpYbc/LUBLxPfv+VE1
yqKdYqi2zhzwWn+MxgLz9pNtATOwvIPPV+jyGTcPWUqXfYDdH+tikncGUK0G/kyndUp75jshVX91
mFPpml4gJswshVCM3hOp05S6gYBrBSu9tuHNLh30BQp+L6fEoMGTMkw43RYNIb7YF8thlTGy8TZj
fS/UKNo6ppLcESndfrG3V7Cp7WwG15zdVTPrx0C6NOSxJB8oUoYOS3/NJE/Jg7QRZxisQ4+usnIX
DxEuxLNqL5/wnD58FHY6KwdDbIlpRKrVTlWaWKoPUvrP8gunUQK2+P51O7pZRs82yJvwPXuU2TDl
TQjTUvwsQ0mtSFjtkkPopGzDmv2N+qBNS8jpDPrTPRLR5g7mANz86vBH5G4kpvWt/+FqF/6n7nu8
RNrCIbAXsbIN5jtjnerZZgjIKDTvzlEFUph6ENdUXkN2MfhonbNF0pbocxLDNJcqukrNaSWkbEIl
uj3vFRzmHqQo4BQjq2w0whCuANwc13u5W7nN8bGtU4aXhYxTSVy1cogfuqxy2P8oRw2xBddTCtpl
ln0hxOOUkj1z2eT2ljdt0g8ZCnMBSKaWSrQIPRxhXtq3+YNVKDepMOevF+Nd8UqyRqavSzp7SN4L
U9xyTmLUXJVoXNSAnZwis7pr7zNa2s8uS5DDClKtmxRJKSOzAgSYnmpn/AMhKNsM56geRWn/v4zd
HlcMpPLvPZRyfy6BdvBPPCRipzQckMnI6r7gYJ4VG3qjS0AV9cnfSWHaFjkoXwhmka9dmZoGzWGK
xQze0unQzfErMoz/8kJ4MOLjzYV67IJ4kI9iOrAKrl6OOL0mcd1AvBIDH3QEjFqYNQ9sghk45Lnh
rWR3cE2+rQyyGyXSTDxQnKS4JzriYMsLCbGd4YijdhVMBwMkJ39WCpivBMeszm1+fed8PzZgbuwf
yeBuirxkFyLd7XOPHv1S8R8X8nJMzGRiMQqHZrG4AaDCdwPTATeBP8wULJuEb/cI9V6EpP2amCj9
RJxbFYGqlekpEyIsDNfzuFcWBoPffi7uPFVH/QgDuolhDhIFab3C+lIhPn1TR03vHJC8BkFVU6iW
zRTI/Bo2JmH5Xp8T9PCw0RxDXeJUSQ4TvyS/YrGusejv76Ettn7LD5+AGhk89JbwTqXgh3snqytn
UwOqE7mXoHvYeYta28sR2v9HepnnPObuhE1ggLYeKaB3qPN16muI7OEjpZg53zpgiZKItSw++6m1
vapqiweyCHiIeMJuXFVHT7E7X3JsGNyt0ZpcF86lnvZ5/Ylu2fQ470I37RRwfVWjd6bLKEiq9HYK
qEpVwzrV1dY1sGCY942EoKtOdaw21rB1nCT9rLog0H3AcmFHVM/svB7rEn+jNqZ2UXj63RdifHgO
Gb5H0zsDBetwfSHgt2D+ty7YZqemC5r5/H3AR0ORtjZTIw7WQIS4bAuGigv01du5v3mz34IghVbe
ePOm7rwWuwfWZv8DJPIybO6lIu2Bmssz0uD6Zj41ZC7J5Ui8+mN00ZKCT/2k1H5Q8Krh9w/tztPu
imoYD6xDlw/8+ApDDUOGpaZI3QN+knZoX2gHNM9V+mjcc0R07eQ5uvfCy0R+pEpJBUlILDouoUoh
yBT5wSfWh/jDEPsbfb+q2iLwSnPr5rfn88hgOrCwfh5ad99/sWIf/HZd+FJGoBpRNaQm3NwNVrz5
fTKsamTAEu/5V2VozjSKmfGULUlDtpe2rw05vWrE4cmU6NXoA0o/oo5lgokcxilUncYtecV6YrZf
9gwrnxMXgqOzQy/zTe+PMi8tPhwLfVpSVyGuYMexi23O0JnnZhpsgSwND4RstFX7prbu0NzmZaU4
tyXzzgT/tOfzPg1hf3M8XM2O1+FU1POgXhqJKLbzhc8mnxJ/cREBP6YuT8wmu0CLc8e1JAlhqXuu
2fR1q+kZlKAANJJ9DKn7FfIp5wpYFf0Dci3LWNvUPuvp1KG8/j/8pz4mrBuAnvuFk4Vn4dWzoWnw
b/6+YtSroaWg4eWOnEP3o387weO7pHi8gz2uW+9b5ID7H6rg5DDvtKTXpAUSXOnmW7mYaH6tZX1p
6j2OCjfpZ0/Dbh2UWYIK8sZlukl0fNekfiSaHCntQbOxX0Xgd1LFYfMw2whW6u1u4QsTui1LKSHM
gfLuxKk0mFqLb1SXHccQefhJ/c5/QStHg83j6+hinAWxxR3Gm+lEdkwT6D9+uESuw9BQRvlFHVqs
XXYeb9/cgrJ7+lIFkvZoWA+rA0pdOWuIYrQGwZaqPjZElkw2G1+aNdXkIw0eDBXxnzPGFq8DAMsg
zQK5/+eSxKLeBhclPNvDbyzfhDIgFQIz5MjYyHapMAfqio/rJhyy7/8oEkBxG12LUxDf+Pvlt7bf
u0jwiLoWR7+mx2qkNdnBoPK7/8xwX9Ao/h1y5nHg9+xQ0QmBbepDgHvQlLKggcBqHZAQW7hwIb8+
L0+PGsJVtQj63NaZ2t+63BLCwZE+Y3/fLiC/a/tUBczcE5KJG2PUAlLlMZE6sTPOIP9IbGFoQkyA
jtdWruQuF5oLD9fAROU2PHDfbE/OKoMBW14TDwkehRDg4sTiEy+MznURI40TUZh9yjOuxyTIRe26
EkK3jUVyCT8xaxwZUziP6TqegxZpNrPGOU6SGvTVV5zJoNh0kBqTaB/TYRhO5UiVTTr7qT7nim+Q
iCB2iucrsPmgEPz2ojIJbuUwwNPYS9XhhODN3UJ3HU2TgP+ixWWcJKBLy0I2oP1pH0oWxvDg6Tip
7hdHEQoWsY+awoBLvHjlmShUx/vkg6qDimT1OlnnCtyqfo2oMQQ0/JmU1NunngkjbW2l2PXc9Mr6
aE1Scv4qH5qHNKt+etY0F3k9/jiLLM5NrWQZaY3DrY50c4bVz1/36IOu/DrzYEkI0x2vrOVBsLek
hRtuUpDfzbCsO5ivNC71D2nKjnj+GyDoGD1U/Kwd8fhKf5RvX9DfA4WN1nKVGnqswg1ZC8sDTlVR
CV0Jz+/AE8xLxe6jW1a/zPMA8FbBEokUe5ShvYgOSlohC5sDWVA5T8W8cX9mcTqiPabUm6Ihy0Ze
iZMnokcVPjwf63o6yC43WcPE/gk3jgWblkGFaHFXkuPwoMY8yVdJT+60QIXymf/fXpWsTXKIBPIq
Kd+LholH4LiiejTRvY9LscvnD4Xe/xSHeHmer5ND1DZg1OJcTj6rBFpQEN0SAek+DIcPmdySLBmN
ulCwd19hi9xDliciH2Nb/kXxVeVy8jg3ced2jrMhm4MkYNz024115FMGR8FBF1QxfKm/Dej7flJM
Y/3BvPLPGaeYkAs9Hqi8hET0vFzebtzMf5Zw8aETI5C8UoGDA5jrb8KcHCIc0tb0rJPjfSEIRt/Z
x2Omz6cvhqHWIhC7Dm6yVkKFjgqneolpMo/ti2UIO/LF6heKcFgU+womYtILLFhb0g11bg4eGO/n
QMC70tHAC+NtHEcwRk80ckRKUIBx/RCB+9I01t/2E0+5b0wmjWOKy128BKr1HSlz73Ob+vz2/QeQ
z1iIz6xw8RMaNfh1HrpIDA58E3RY03sX38Lpwdj1cIz7hwgFN6QxdZUDxLjId4J3xlTGMAkSq+eV
6jgYfk+YCG7tZIw8kKAgcjKw/NEtaLZKQC/SGKhtc/+axrbjWKDgHxF0b+rOw7xTJ7Gn8OGTj+Kq
F9LXMPAAPo/MSGUgRRn6XnYFTUMVC2a3ZZ8KL2mDUv3Hef5Bu4aIyMNMYlGYN4PPBILRyQAXs1cg
8BvECqKz0T1FqKzPbJyEP3VOnNyamn5EDEyuXqZG4h8N68EQcLyahZQ/IBmQ8eAk0zVlweYc4fTt
3Aw/8hwlcQ+yxMVVom1gDENXwEwGrY5Sxh4CxbyHCd+inPSUYW2MCBJQjCa1cUuKkf7kFAu6+b1G
blvmLMLmLOrjb5RlCgY1vs94snoaFUfaA/Dwj1ZMVeiDagt8B1tdjRDOaPrz/nVIcx9P5bLeQprU
sxdlDG1hVEQqW/oZI49YDhBj8P/2vqsQgjFTnG7FHDpPWjfriUXreXKi55KK4LEg2uQJFK3BSSYL
7KIikRTAOcdiUQXv9n0R4I6xXujrVOUmtkFm8Y1wn9UmT7WwBKdyo7NO7yiiNclor3HVO9OmH3tN
SxZ2E+1TEe4bdRZUY7I5MOMjppXHvjBtEnlNUPUDiWnALiwT8Stp29oYlxWAowOwhr7OTFu8KSNz
K360juWKTEQ477mAdVtXcyu67IhBmCl8L1kTf7OQlssJ/+RrRpAK+/rvp6b3ILdjroZ8nAGq48iQ
fh3dfdVj8bpqhycDGZMzXBRxZsdxRbYJ/C9zWLkBuF/VIfvZy1wy6VTCExr5riEuBENQWorirurk
GLLFE9tvtAgEdHbbbgL1AGoPnMHNOrS8TeSR9n7RsGXQMQQoYiZAXK1Vh68wp8Vpc1njtpv5583T
geKgd0xsoeZMvPfMSJgBicKcMSbq3An2pJTAgklQtPdY3U3EtF+JwNq5zT24xr0TXMEJJcE+a4fD
BN5GO7X9Q5p0F+J44FRBwpuY5SnYSpQGsoh3Nq83qOwkVzZ1d/3RTUsiAUWusQwG31RWvvLcV0Pi
/w8Swz4qLG+oFPh7xMStDI2odjKM7+o2l27n6Yio6jpqE7lCUhr+UnUoO22yAuZABEGFSMDlz6ar
sd92MNkPdjcdOCB5NFue0gBaLlXWFLBydr0xq7jbhZgkGBM5Q51t/xhOaiOocAWNyHqSXtaJzny3
stcWe2oa4wb+KmdQw8Hf96zefSbBlo2uIBuEREPeFixRi8RgyR713i/UrfnrnCaDz2XWi3143D9v
UD1treX663iAmQRwpqU4X8ZUUp+y3NMsnu0L1kQuu7mOA4/UDQ0D61zoZtIzrGgbL5blcpgKdz43
RqQkkNRPiAiW2tbEwW2kIURyqO5PIEbHXXZRogVV6cLTiY9sdUbJGvUiQGRJwT2JDzFnnBbZBB9r
Zvx8G6V3Ndllu4R+xVvih73N0C3j+hOCv2UwO6D/ZI7D3oQd3HsMEYHz3/pERuB2oOpq8JdlNh6B
AaFrsV/ksgXH1r+KIVoXG/4/RlAI1NUZ38JPyoX0VyfDDw1L48hx7D6v5KKn2akITUR0U5B/GKKh
2KQchssJXOQK0JE96NNZXYke0i0NIzBVSWBobts4s/hJY/+kEV8dICU9mjUqDjHclA+86JpZpcEh
wKwkMojRv7WbUN9rZidf8TdLc4NmWh0o5gC3l5cXUdb9NojheenZ3xPcv3mtM2Bvz1Y5D91hGKCq
HLoOuixq86S6f2dx+T7n9dbgPwVmgSPjqhZ3wK1vIUw9cLto3G49uIfKc2apP535f1MZYXt4FeMa
bi28lOmjvlxCt9SbzTd5TVnj4yr0JAEl22RtepBfPI9o1h65dwCQglx0ac3gylbOJ6EAP9xelN/H
Sc/oZqTsrQKBJrw7KxFSM0ciY5qT47iIdY6Dno3OgRoQwa6ARbqS1fMZLMg440dTi3M3se72A74u
pku/qV9HLLF7SeOxxgCUMQ8iUPz7RHbGixkDOTZwhvMgxn3/4r1mJOUzfTn9SDBl/cpGzWBesfoY
/yiH9eJ+gdDJ6q2lZZAqtEBBVQg0CT2uS7xaFeMGUaZ1bnQ/jiJRY28sxD0xPOmPgTv2VXayPRTS
KRgljfXo5LMHe3TtHO5DNr8Le+kpjfnD8sQ6XYHSq/B65mihj2J7oXR0tt6xx6EeyfoekEWHqCaQ
KeAsoAwkS375B+SOpNxp/sMLW694+F3PyMSIfoQTtNpfTmkMmsD3nncm7y/ZED4KMtvyEAZ1JupO
Or81FCvbBFFqfbF3R3yTdFY058xxF3Lit+HA/QJPXQov7Izh1OCsNwSRyL7NC/5evCbhxnV27qtu
hSxZwA1TGo9IkDl92FHpGcNVl6R1WB0u38a+/sbmK6PgIc4uC8y/SCrNFZPXatnRJUpoR5NeLnC6
nZuPWggh9UMkTMdKY/TVTqfcivDQp12x9ygn8tggaHj6P/FybHh0q05o0TkU6z+DyXXp1sCgygeS
a5uK8WNMH8axD558atdfTIN5dqWbMnbjGH2AcdYuo8vKewsttYuJu752ET0GkFb5tEjHOPkU1uyE
+J018gpsU97UzfdbZjUvqyTTCbLTL0iVrpzbuU5Rxnyp7AutHF/pQVUYy6BWCrOibxV2nVV2twbC
7a4C8q7zNoe1NST3AehX4UzR3l3qUqGC3pEdfOBgeU0OloBAEmtAVXjKHiUDcgzKif2emtq+S0fZ
bpxNJEyhwRBfpr3ZWxDfrhP98h9BX96NRrEJFcPI2NxURjPopYXUfjPZZwPH9gUCmdKmZNP/FO10
c+TOj4LS6yU5uD4n1g5zPm+rzct2ErGyIZzoxXY8ANFnoNMy9y94skasAa/VdwuEiehiLIRsJ2f6
S/ZgkgvpudsnrUJfISYmvYLXX5RLdbJrAq3t5JUupYo5vETwgFvsw51IsgoIQ/MtGF5A3qOpTxUg
VO2R9bQMxfoWd04dh3niyCWtDQHZUC0bqCAP6h3trzLmFD4zyc1p++CJZat+CnHziUz3f31YLWBx
k8iO+r4C9NZNOx9xziua0nSM6XqmdzvNYGNbWxrtPvae7ntwnP2juvRR4qaOCW0PAy4LwxvrozVi
ywABHEnYbG1NO1hfS3yp4UaMYJ28YREOKcbHmuTN6m2Rb0zk6S/kxQTHae7hiMaYZnn2nCIDaM+H
Eq7A9GjpajkNVFgFRuiq2xyPQx9nVbtdOicRx8/5VUYjvY9yTKv8WoPLOoNnbFDtjykK0wxa7OAH
imshEbqqyRL0dVY6zhcjmYl1bGTohELbDAldP6D9ptp4FsbXUWP8sqedKgkyqECQGP/N2xJkAPeM
nH1CTNU7oi+a4jArSuuAHK70QhyF+0Jz9fn0kN/Ft3KgUraoWlHsnfcsGBl8gWkQR8+JjR9YvVgk
0Og8ez97wSBKJ9H+5F9XYCFKYAnFBbDDZoMTNweKZt0rdIhM+Hj+FPqqZ2FCxedzorxM0NNS5F4z
JnEz3IGQk30AUN7zLujXd2qgFBk5nSb2L6HZSwUAIMmhX7g+uhHDInUJNVxJ0fLJ7B+lSij2S11J
JCBuYpL1upePeuCFFJrIrx6nr58d2y3hf+Mnfqx7PBFsECvJpbJ4bzdT/cDzKInJ8oYMDyihDBaS
FtjMCRZD/0vDlD2kUIS508dtdhhD6teP/q6HOecvP/6ZQUL5sXzhhTpHd27/GaXLmZQHfkDqOHl+
n/4RWOFm2zzHC32emK1o8eZxPxTLwmITHnYZR1i6U6662XXqC2RLT9/N2sw5WGzuYXDViktqqnBF
WoSbirfrKnm+pYvvuc5S19ydGg1QmssX1QcIQGbpvknr3CbXqACEQxBsO4726TAQOlrPiOQ03kQi
igXZ/eWXbgzlVs08MkKwwYtLGHCGSxcAvNjPcVjB8Qm7DOdSJwVlMav7dLTqAzA4hhGpTkEulNHT
FvNrGc2uNdAjocpfCr7y2+xGHTucCSUVNHDw1OeHyJxlbZqsdbtR+pVsyfFyhyKS87Hd60VNIHC9
HfO4Mv8ycJrYykh/6aevsIOe/Go3rNGvWQPs0m3iHTBn2CD0fyGjvG2GSuMw0uXLBtIPvz3+NCyM
sib0G/TSdcd4W9Jut3UZ+UcYJrUWEE5nL3JHQueTBEQL7AxJ1rRCtADf3JYaXCsBGFjpKsW5ctkO
Zu7AYZLQ/c9GdKRl9YfZp35fiI9k7K4gR2voetGPLFlC78+oFYeKHFQGSQGfGQySJPDtbhSzifal
0czEnyhi/Jp8aql3ZE3G0p9wmpuqaqm28TDvv9RCt78sd07QwYgxnwEo9fufbM7jy7djupHfYdgm
7RHJfKOtIHCl662gSnpgqlkf0Ft6JXPJ69wFspftl/GJNxw6l+cyD5BS6F5CbSacoMJjrgDfpaQA
6KXeJGiMi9j/SdXjN2p5fuCwML6K8tFBLKdyIUn2mYHRAzNgYklXy/aP2VPFID6wMoaiZVc5tGw2
UqSebpi2D1q60SREorPE9Q91obSM4nSapcxccR8y/F7nJcCGdi9FPAL0OJFNOaAYsUvN2txQCWMU
Xo4zaIQcUH0+Z6CQVbNV7e2JqK/m90z0JgRn3i/vcbAfIT0uv+Thq7KzcewUsh65MFSCIqu7MgQ8
F7aVs3Nf1Ymqaorrwd5tuHfDYw8bpvrOwkICIenkp0B8pZcAQrGFZNTeAjVAKlDA68vmsbRNRuAc
jfmCpcsvTf16T8sC6MiEQfCSRZ0FrcpGbudE3xeTEMSDNLO7QzIA9IMeQkyw7aY3OEuGvZQ5HbF+
3mf55nrQCi4urh4x8Wk9C55J94NbuGOANhDPX/KeiUoAzIQ7/64tkx9jX6nfaM4bFDlbeK+8TNX7
mBqHYEVC4oG33LRxaaZgs61DaNPHoh7ltSj5JbX0oGBM71sRCuElnk+73dXMH/MZgRHEUoddtU8a
XPOwUFIvmuZ0z9UGjfBOcfmFeHQlNwxpxsgkQWTjFwzOSmu36RVkyOpcwE1I3iWujVpt5Hl7DzEW
oCyEtmjVXJe/SOSTQeEQKyIcl+plVatN3ZF3kB6mJhbVAVx/fiV7mUbzgoCPrrTi4YmVHcOnd++v
5AZ5EQp6WH8qge5R8e+EvYKEu+pFv7gt0vEIEBpJ9D4MBZl4ItfYXUdrwFfqDp07XNFlvU58lYp7
idDyuD38oM/ul6x+NJMG8qdrZDs02sJCe85kybGBaBoW1UC9aamfk+i6+J/ku+dbPd7/OhnweX+m
53QHYO081HQRYz0eYbltwVLezWlD4K+4UiMpqy6Nl1XIfK22CGlpg7IPGxYadK49tNyoUsWyKOyd
l9SuMsZNTD7qfeRuJvzZj10ZZHckUfHuzNGOrA777V78NIPqF1VEhU/lAFu4nY5PZ0ZEgOU/IYRz
Y0pDFN5d4GLuI+nPTjxvkx5kLgOc+BNFyVKX/WI2hooSBx6UCWsT6I0zjTGNH4YJsLHouxzX6I90
L86N9laq/puAB6Q/K5UGmmVbqtpl511jmatlJE5J1+p0BNeJK2emMpfwrihQeG34qnoKgnmapWLj
RMI90Y5vTBLStNyx193M1huwL5e9FzlE/BvkLVisAKsIiU7hPNzoW+CbVdgMGnrEDqMQHWSj41S4
8HuTeJPwoCsKcGY6NV/kNWwo60SAqhXes5H7+OSn/MZT3cnxVQgGMXWdH7n+l4LyCRhe8ZuI3PCg
0/vZa5imldGxp+WeWvN24k9b7OU5lh9kRirSwpwwviV3BC5p6Jjhb8tSRmGTKQsQmN1n3UMUXA/D
B0wn/C8r/wiHxtsRQrw3pFF54o7hvKUZKtmhgJ3RQM7ypDjrJvU30gUHI9NnsIvvDBY1o6I7NrnC
6FfwljXnxpMfZfCWH4FCAZOIIMl+r4MAachzr9G5F4/KVW0kvhVik7tcZ2aY4H5YR2UugLlrkpXo
eMGHq5XPQIWWVhd0Zxly6mm48g9FrGm98Z4BUvSvObcyJ3ktk5dvcI+7a27pQV8DLcfS0R0WxR5L
lF+qbeGNPpXcunXD4EDmFkHi+qidChR2Zt2YfdozHoQLVDOgNFFSd7BgYdjEOSlJh0OerHoYyl2D
ap80rScd6bSHPJFoE4ALD9kt/a6xofVyYtegMZUh9TuEbEQM5NEBh4ooixgOiycvbplPcPjcT/0I
yi9zl9FElIucFtOoJ0fFewAENPkS9WtLfcNMoKtCnpFbo3EtBwPe1IujADExX2yxXs6lefpGp99U
ZLt2C9Dw1SL+GJ5EaT3aMic422FtpnicKMrFnBqiAS5oyLzFX9PQlnw+ruN0LxhHQCmB7CUseoPU
Lhr9CtGOvcpsrAsWCHn3EYbxjG5tpqWsJNV7x6wGgL8UbFglkUts6L61NS7MFIYvKIXW1ukZ8uqn
JRxF50bMxPtmnUGwydtvWAARTp+nW2UEhmAN/KYaMf+i76CGgVC2oxosxmZq3o8f8DSBDDWkUu1o
H8QtoOkUrDHp/uynaHOofyvWh5AmJbzsIhbckFo71EZJpCqxd8Jg7CDXwDMOqxPgawQiRAnDkGzS
zEQgS61QTnEpm4tSRd3Z/5uiFngs2dKJFSmkxiCOfVJhGt1WKwIbWGZE3YjbBm9chvT7tzZfzp3s
3ZQgj510PDmbP6uHLZm1xwAZzhDip95n/pXco6MjLxyKMDGs5W+ymVJMBuozcO/CuTh8xPxruoEz
V6qIXYxmS3jYdKe3OF7zYlEww3iXaMfqkYLwdAUgSMVXEzzEZ8Hb+6fg+NNVbO/CpnElIo9cf1dZ
+xXqOUbJoNMydvrOs49SID4S23KjavmeMaanlj9wEpd9LIC70yGbyY2QtQjFqOhTd1qmpRgqbCGT
QEEXjcFqKBaI17ZX9AU34LVPoeDn90xypRJDgd3MlE7J3u5uxuM+QnPSTtngp4gcWOBcZtom5e7Z
iiK7SUxdJvNnsw81DN82VyaCZX/zK3E/IpzR/Bg0mopVF5n/LXNQccULpiBEaReK0a+LrqXeDUyE
E0ROdMi9agsQ8+JAGda2i8/a0s6Y5F+uNfYVYTvOp3u/QhhyCX+EZI8foP+G6XoCC1yEWx7YRIX+
5FEDcXA5iYzC39DHmrZzjE7/oToemGrM9HJCUm+hX+sr4jizS+3tdM62rV4eL27bx/M3jlPUVXIk
PvQ3pV24wOIJDOaFjwbqnNsMMeLiq+BG4311ncHq7IHzDUz88bvG0OUoYfg4ZtcdFNGA6hElA2dl
pXN2x9qG0J8uwBh5pag1bcP3ERdW5dHXuOMqGJXM15ns/FlIxg2yJTysntMh8GBqMed40nFHFhAF
koTv8dnsqebV25kNgbHwGuk/i+CBkoWQNu1hyCBCgBflrQ+A1Zoc/yi9cjteUYFK+0nB3tGcB9gn
BCI316nmCImGiRbD65epyR7uZwMKCcbUKG0LClG19eQGQf4FHyy6H1nHb58IE5EIZXj+hqblv/jN
u7XIYsqng6JaFAP7Io9+tL66eaVmkTzjtUjcLzg4+R+m9zoWZ33q1c8u8qpykRwHoFV7EYjiS2Zz
ueaoY921Wj9YQW3TXfv7AJLvFMqj8yFbl2IGjEdynI4f6UbqthkETHlcpvpUN8W00HbbxOag+skD
ATCyivqJCHSfjE0cqrn111sQ97X3hGTr/ofU6/RJnsI0ZsnjoYGiVDTo8QymnlwHQ9uVIlW8KHOt
nG4NrAev+gwX+TNqGIslZGhaUgPvayLoePCJjGSPuXxM3LAY7O52sudZAjjlc46atWZkxnLR6uwm
YI7xdlfTNo4dRbumjPKgTStadzjm+ioH61/EV3J61Bz+uIR9d9gWihyHlmk6Zk/adGF+lU/Ms2sr
1dQf1/4A5nSvL5KWn5E8Y1JLd/iPP0hzpSiK9CR2Yqh+5rAvdwbaJupvPUVObxAdvJl1+X0IekZp
amcUSyf4/o6ytqQxE60c4FFmbnqz+m9QvwjnyJPf6JiBWu/wvQCU7+LogeshhYvptIRUcVscrH7V
OkKjJme8hSyzIgt9fStaaIWwUI9ibI3RjtWHjAqlHlnslJf4YGIbORfdOHQNKCuPn2ili4HLb4BM
9HohTXHWiTip3K1eb6aFQkv/zH1vc1HGHcPTAg7OPkt3Ob02Jqfxv4eT9RyPllXI+BV1FEezEUTC
aZkuA7BhgjsHP8Xgr8R3c8xVOHWCuh1gIOCUvq34oNwTv01VRMybgTv6BuIelAachsDmMCEIiWS7
x5QHmJ24Ab4Bfo/Juoo+MPsy2Q3/UgHGNr8L7oI9ks8QeuN5aBO1eSZwFdxSpSMsj+AFLgiEzZue
UhVOrYwShv3jEBfUm3hqL2pNwznkrKQ+5knIh+HeKI0eI4Qy6OftbMHlGqQMvX3b9TC+MqRlU5yF
7ihMti3n45zcgSafTznVH2SdgoOX83kCGp2L4EWsD+0J0d6sY8fs1hbqXRIysglj8fU9i7nEY+ck
DGdX05hpdez1grJSp6V2KcTYhQs4P+ds419qp+vehteLMfaTIUeW4byS7fIHNmOdzoL2kkTg7/p3
JgVs0dvrUPhiu4Z/uYK6eIFssDGIuiPSdQFPDbc1XgF5yrY8oSfF6iMtyly3RebO+yMq7Bhus4Fm
jmLCF92mqk0VeYWEAHkFYrb/fkGpFno9DyTJFzMGi8NA4bag8YcpS3ebUVrNDv0W0QFqjw3oAIto
XqUBcnF0UTZw/nVsOsg7L81QVQfXEy/da7RfNBFQd10OEU379VVr+TFKednRykthE/IvbA0LS7zp
MUYBt6yKla+l1TEE5KpL3dR5O8uo59yktREYUTn2AkrgIHARMJkOdEhSlGuT1I1Pb5brec7dJfqt
pMplErdPLZ/4odMpHw3PVHWGgSpSTxCbmcoabkVJFooo0Vdha+LdcvY/it26SF9f+q+XbYf8PNyt
fZR5RQf/82cTBBWFbRVXMVWBOm0MsTwJPCvvckfISiLSi9SAn6RRa3/ULCvVxhadBhUQliM/WOnr
nV/H7jHDQmzdsM5ytYzNgE9vAvvxtFUnpxPMoZj2kRAeH17XYo8Qoy+syLRKqi6jhCKxcQdDXY4L
DVGAVmynMtWzCmcd7N8zqhTjpNFoGnfV70UW1X4YGg3nxeRWYneqcBK3udZw2DgJnYgT4rKnMxV4
0EnFFQpnHnNhOfC4Lm4nP2LXRP7OwmSf812v1TOLRrVP7aJKX139UBwQxLBoaRdpVlRj01QMkqLS
IPkMMVI0Y9ODMCUuhSAZYmncFAGfjXr8kmtH4PZ9ugs7P0lJ1+TeouVsPkminUv3GNOA/pcHA/3q
0GVWaZPOfNunXTvcohXfXA/bEM30kYX5hAw2ht0Klx9eJn4xndaEFzIxhrvZv1il/K0tG1KZJhFs
aZNGfSRrp0k+pLsKF/apARU+djg+uA9cLoow70xbvDVwDDWQlbhDfcb4LV2ASJmGZUgSE0slAuPL
SZtB+gRKrrn6ChNMoI1wAHpzKevfViTlCqjxCyGCRV/Q2IqszYlF1OZDA7dsg45mFKAtaBoEEd2C
cy8fNdqZXfaBWRioChc/0o0HR/sbKhhQ4QjZ6wJ3RPbbA8S6IH1Nb8i1f5+sLe7OcsHGPlYSAoOA
sVbGUlySfKlsqMgqv4cdYIRZ6XS8jJVOw885QbJAr+QclPrj9tT6Uk1+eF6FpyGUoLlGEHFyTh/X
9kyodofKVm0b49JcSwHEpxHXW/lISAsGIUxDbcQVFHS9/2KlNx1hI4YlL0i1ECmX5mwb4u4mPocQ
7Hus7d8A/WVz/6a1zCumvec1LnMUQA2PunnikeK0zkUnFF7jEHn4bxdxNOJfJsuW4p4qbyRo/owD
TYDuSrnIo48N/o2TQ8s1ZZozblpifGeNg08kJ9JE9IU6BTACCvkGsnLnGM90Cvmr3n/zPUSJ7CVG
32AResyv/B0o/1XhYoVAdi23TPM4rT22q1sofUitZVKhF2xZMJDhVr8yS1eEe3Qpw9u6Isj1WIKO
6u8hAEouUMOgBeeYm+Cnc1kCmTjd/Ip7SZsUPUGaQ3akY84hFXlUXNnUEjy6Cflg0FfnkaTUN/RR
HlMDGdOS8P1htgg7NTwt5BFX82YaTC/5pUfb2NBbNVAtnTuACaxVr4jnpzuBlaMZYuWCPy4MxELB
NQnor7Irncp1B8ewIGxZOWQb71bBe9M8QMibdf8KOMJLHG86syj0yMlbxkgJbo125X19TOIa3ZRb
f0KcganzRk5BoLiuWyjxfSyT4+bFhnYZ3NMuyYzZ1xEO4yt5oA8mGjeSQSl+F9qpFttOvOSBWZKy
jrfad0jNALpJ7RCw+EjnUj66UxPvRp3+EppADPJiSOfB3Gp9/V2kbSAdcjVoQ2zEfJLc+6n1K9mX
UqWruD8gswOYT+36IBd1LTs57P2UvtB8oHNuZc2hm79lEF8fgxdbgW5uPyn+/rSn9GtRhIGLW/Rf
bEIRHJbsXLsFldwaHf1fcGWSNqv9Fa9r2kC/myMOf+fer3qx2wQsQuxvHbXt2R28kQaU66lGuoUj
w1pCKA1/bhzl7XnvcOyB11gih7BI5lCyBRGXYDW/YbA4PQCfRdWkVuPsYej61XIab4N8TBU1Htv1
qmlUH0A/u8hXJVHcS5B9VZjtGbvVMF8vvZplU+HCtTIueRuam4+bcI1Ydn5P096cs1RS8a3SQbaR
ipxuNcHzAvNhyl024Qj9OB6DAxLucgu0l5KJKyU6PaLKYp2Sc7uatC6qPXagnhxhBOeMfio2sxp3
KxHabnaA8gNPGApvGabOi9vqr1A7uw1r7agSSsfjjeqkbvADH+VizMAnn8lKWoHumQ5XWHwMdfcj
TjMOU/btWHZ7B26Ikc2+ZtgPHujJNqXAdwmRgvDEXmHDdvzM4349KmlKwKVZh1Gt4xYKn5e831+h
FrQSpSJofWZEzx6kDrLtOFXWKLJPcYELIrnfWsYduZymnXeezpKpFtG0FE5s/7iWB49wo7zH1SSg
i9jWA6HHP8ELz/ihIgGJ8zQqdQXh9bp3WiHhiMH7wKNDW5ZfikYPDB7hsCqxu+nUQRx9TCYYMrvF
5EpgJsFiBHdJqK1RWF+rBitSIKf1o6pcEn6ahzgmrmyURqYNOfAYQBxnVv+DO6iViKvoxIxqwmEK
yx5LTZgUXoURpYGoNEcqFgBi/x6o3wXoIEuh70yN71/iOGFUfEpYW+goHK9h/1K8fyetB79PUZlL
GzIKWMqVHIL04clhGP0HYmcTf7AgxUjPu8v7mMVaw3JPJsE9qPxTTBQG8Ma9krStiJVAdxAH4fh+
6JYkQti3rPLRPzdDmhESldM4le8NdJkfos5gz6SN+wDbIYh9rTG4MYkX2UfP9P7V9YJZTG3EZ46p
lTvx/morLd+On+dpQ1UJXdi8DJI/TIntwiDoF99D9ritn4MBsfobnHyX9L2WwuXFNDZXvoo9OBA7
RTLbG0yxJ7h7xYwQq8k59HiJ8GEFdyD6ZB3XTC29cVgrI+koArBuKO96YJ86ZoiGths9SLNsb6Av
2xx3kvK2XT4ty3E37dVUGnBwCm+9yKvp0jmYCliYC382EfK0ksAtfKsR0Qsfk7YfD3BD1dsbEFS1
7iIGHtWNcD5poV07kgoG1GBcI0GIsdl4yqm+4yksi/y3z7oRj5a1AiYRuCgchhDBbsPvrjDzprEK
WJdQe3WHttBiQ2l2WZAK80XJ/pVv9nyGbLqtnIRo4XjkELJzab/qfP3AZm8JqrVMLt+a/VX5v/M3
y2gAgH9nYCLypax5VFpBSrHSNkG5q026Kr8MF1Dh1HQLFPnKnywYvS2amZTCa0te85okUatnjqyG
gN+qbnFbMZLTjU9yTgaaUFE89c9e6mnrhykxPCIRchzD29vehWQbj3y5cbUe7Zhl9lkB41/vZAO8
R1lXiyjoovxB329FWLuza+VyBMds6+IG2TFLsqXToeTJ7VZK8wAhxyDa0UJFDWk2Am6rQD4frlcL
HAPKEsb3crPtkL+3W5//V1ixURSGa1+4q9erfk8RZBo9JZ030aWm8QvtbvmOyvhVVkwYCa7aNl8+
Ch32CeWcbNClAxewRLWF7o/n9969R7u3mupghZD+FLSwtxiSUEiAs+APDJanjvsKBvY+79XUB1Vm
3gQ13GorCuqrYxH2HTONgjRAQjXPQ+yDzawRMo49/lk5J2e2C0CAvgLiAC5FCYCLD9ymhyDzqCm1
mZIybVqXfZk0KbSfAXUACT/1LYj9+1LpUTq/r117V1sukLGbeh5j5joBPFxMj0P9/qWfc3oOqUU4
Hs5YDYhmsS6rG7UtPa8odr0sZIiBT6pVTzHnRBjf9WPTKnbtRmn21vhADX5X245eAPOqPFRELIET
jTsyvEe9VQzCJbYSaqSPiiGGRpqPIgHJQ1j6h8AyJq3B4CUAD9N7/xLLXH3yCWfPUk8Rrako5mji
eqN2EEZ+pVIv1P1oJxymoC/KLNvq0EFLyBdDIHZ3ogauLtJrz4upCSyWhPs4Um0vSsFHqAB9GOqT
B3PYvmErUNbikMQwoUwlyjvQXdm4yZez+4Jh++xbnJ62vEOae/y8/Gzhly62hxSPD3/lkwLQKaBZ
FkspmZqKQXUhBiB4/yDuLCL/JI5EYTdRwWRbJVMMyfailVpdzCwY7YUvol83spzQKuaTndfwaaoX
chDyOY7Epnu7QStxbRpw7qsU2n+Rycoge9DPaKDTywZ4a1qSdYSgyE9VVtmTnjYxmiVP2nMlxJeZ
TxMh7LwojKDa755xqcmrYcxWk50Qn3dx+suoi4oO8yb8OC+s8l521IQY6rLrXosVo5hR2x3bUP4T
GsuWaB0qJW9E0m7pk2s4UQ/yL6XKrkqJMw01CYgtJDegT6Nhgotk0++ah6Cb1sVD1f+UEn46icUn
hn3l7ixs3VyZFx5frgtf/EP3p4pRXX2gtcYgscwDLM8YiFATcCXrfEO6itYyiNg3PveMaLsCKpWG
Mlh45PAmxjYi4OQL5yd5h2Zqz2HDdVkh9vmlEojp3yK4mFumgfGAtoRIzZctFmeaksvQE5UeCDPD
e/Xb2HEkw+wC0r+MHoLYkfrbjMqYMBJOtVUqagEc1sZZwuy3wRI0v6x14Q6ctsZtgTmA1yBWN14B
Zn6j/TidP91sPbgyLqi0y7Dj4o8rpgKzYfrMKr1pfaXFohLaFTGZ6mixJ/X6aK3B/euLCeHwxzpE
BKPmaF/JGZZR8LJIj/1D/dkg5OMPB4iYk0Fze0IVDN4/d5FkS6LIOboV7lr0CpDO76Z6q2HHzPHd
a6HHMhHn7lUxC9ejGX/zMjzZ/NWb2xqbo5N+XtcQqnsHBdUGvrBfyxMNhzkB+F80XjdiGdQumelQ
I9cF0ksYHkys8W+myuPQHEwucJjdXnW7o9ucWz+YfycY2RDdsFtmZ6vuG3O9E5ZWYJNsFOMlgIeK
aPYFIAWYj46utWyax+lYUL9S0xZOMJQQKGEffpI/K3wjBj5qP5zPe9+3HwFmgS2fPv219b5J6xoB
qPXSwnfqblvSELIQg76pHWc1u/61NH4yxmmM7y8cfFrAJe8jiXcOGMwnaDw+2uHv8oOlcyMdeO2t
n2kNvG9kJALa6C9t0F1Q4iK4J5KdAYronwy9f7H6UmZfmqLTVz0t1gfPyQllxdvhIKKHSizA/D0J
5I3g0ZQ1cj5fEtJbiW/Sknc6JY1ZHlGt33eidJxv7pGAoKekwHI5bcqc/hXLkJW4VjdeE1VZzwCe
ds/OY/1IA1gEaQJmX41SOl9e3B8JDMUXkOy2xppDvHEW9c++3NlOXpUUql7lQpHHjz1W23atv7nV
eokzd+LBUF8uaYneGImfOScAvLMIpB+c7WTWuRuPeR9fSHnDNZMa5dIYIDrFS8LErK4W7j/X3dNR
BbNAcJ4Crq1b3rGwpDIUiNgEegjbfu/52Ikxnuh187dM27pm+aPeMQDxPeNbyd9ATXpBRIHGxv2P
plbC2ckwgCtVn1gPmqXzXgwAlHhVbEgq1ZkBZpsXfsDswCq1AmR8eafFJ8BkFVZ82f5l5NWSf/2F
7mhuv6/XzmJFPzLjkDv0TD8FzoyUOTQW/OIbEX5ZLTZCI9BzgBcU/yPy1EyZ55rq0XVSYWQWtm4a
uCp8uHK9feK0E3qZdJiJ+PmCyMVTHFkqvutkQL68s+OHGQIeNTCqXtQfdB3Be73NyDmIZUBSfF67
4DArRgs3DSB2aKPYdJL3rfNxsk7+hpeVvngfjrrL8Ex8y93Z9Qz1fuFdglD58/s7RNhDbeCxZU0X
82sMc5WO7rtEcrlmJNK6uPCyJceAjvrAiU6bTH1nqVWi3kzwP3roCtq3cs+P3iBghSiLE8OTZeme
N30fX2Jftsu4xO0yFq6NUHKptq2azYS0tslFXQrOYIVTJh+cXFJeND3iQSdfyJb+oIFrzyLEfCzm
rTD9NUaEu7oR8KsawQYpBPNGWnMoqeVBWMBmagmImbg1M2bOXicXok4go6bnUZsORLqNOArfrcF0
c2b0RaEmQAr3b7fgsJOvQpD5obOQ7rtnnPgRkeEEjDMa7VwRrpImdScEmhUQNksNqDzl5Du7sJ7k
HrM/YSsSinBB+BQBfLXfxxZCFZk21AxuTDU4tQOPQwj+TfoT02EdGE9HYjpwakdM14h0S1NKnoH+
lJVslsLaccluo8uyRy5u0mcNyJYX5xQOu6Zzm4fJfPVCDLu3z+YRpkiWt05yoe8e4UBHG/Yf3ihC
iAN7+L5hjBCG86XdoGRR/k2WRu/CWpamseV0xlX+4fsKFfBSsBo1BrAnUkWBdnpntUP+OsPsWAz7
XIudYuA2+Ix77sMllSgEFrnFWke3SmtwaLfeazIjxO+WSNYwAUKYLhRSx8QLZ+ZSCDwtJV4qclFU
G45QosAPqqExB9KHBoNEq0UU1Pdax2bx47TPg6c1xFg2rBcMmpL3O2tAyXpKh54ZFLwsFuJV8IYG
+llZMqiKtypC0O93P4AvVv8S8eB9bqXLCRz8K23wlfqcgrQptmTXTaRWWKkbgE+gOl2R30NtvTxK
BdCg+dVrr2AUppXRGzhngwvp8ILm/7G4zSwZMA4eP5Bvf8nhcVWv5NSXELGA6KzP3T1zr3s2n9ay
+vr4JG3hwokCENySPqdou1dEGge0nOeA4jeFD3kP30OCDdtdo8QScPvFI6UIRnUJhTaxaWGrmfOY
TY3zGIh/N3YjFiPTiG+tuMgilwYTIfhhf7/plguw35XfUCUkpqb9X5EEJRBTODq6ow2ueC4zujM6
EETUP4stRUcHDfV0y0nNTicj0uywK2IWNpTt07jLAaNqKhc6uXBic7+3PwkkoctFNCijTd0xZTnR
XMM3I+eBwQw3TLQbZqdHV9cnb6MTo8YZcBX/jElYirM7BWA7EgyYcGJ0hHBGv9d2YLbCwB3iFmeQ
4GBkY6e8ICV5HYnctZWlkNJLU6JB8OcfSvhjbvIOpZjNwqhYlTf0HrCHHCy616+7inGMRUIrJYCd
pc4WZ/pABh0VuJL4/qKU+ptlFiMglFa4fP6z/jQHwWIkIYGHkbwvtR4UwtbBwVyGWuXu9rvi3vaQ
QhddlAlFYkIzhInwrac+cIJowsDX685r7JlzgyPpwRz6OWUttw0lhrVTfN2vE1ppCzhWT0ZGRpja
u0bbWFzS1fSsNeFl66jtdid9uJBXOHEugSUhf0MGkQJvu4suu3srGAy+Z37rLbD6Ee4ndUrUjKtc
8BcH86dN76H3LPiWdXTXEVQMjdCtg58GwYHFUUotspZHfr+gyOVHrguE0appLPwXBa0jPTIhhMFx
vOcV78oOc5c8LP4WPvU72LVVq2iYH8LAbn5P8Hq+zOw0Gq//A5LWcRsdOGwzU/Jo6BCJ6tMyKbCf
Eg28mnTAAMeJoul8t12ATG/GsZSYuLTw0d1IhcHkZj5YCqrXW4S7XBqkkdTo/Q3+g3Wj9nvVWyNe
Z7MwY2lMtYorknXkYPfU8Tv9sqaY/JwCdua23byLv3nLbhcB2B8wmzazECUJAshdOW6LUbtLar25
Iu6VVcWy97Gk+FkjI+AYBiIGTUlDgsbLaS9aQNwCdDfgDdl/siEp+p28/x1+fZwUH7whlEkZ0hyQ
N8mBagfltST8GXnvIc5qTV8ZV5jp2ju48UEz4scGMKAg2j/YFLtyV5C0uqEBk0bc6p8Su8uXfAuq
4gw2ksy6/D75Tbh28drHP4A4IBYiA5QbWOBvnF3UjhSOV89ZxQF8yOZlRKtpSG4ilu0GRtpe/2rw
ZO1XLOig9W3Bgxo75zIX5x8L5l4GrtQOUTMJV8l893GebA2Is18l8Y8DN4m+o5WAb5qLuEddBiNh
y4sJXrZFXEak+EBohaJZ0sqWCK4b/5D0zFfcoiQxAqzDNhkgdV3Om6DBtFuj/ledf/W0nZfzWIHQ
4fnMdLxRpaQUfS12LRJ7rHL8mUt1DM+jCIRVNa92CovK0dpDBTWuYRHs0IRfu+fsVqALIqpSh7gv
JmUIbNJASqDFK12c+GEID5plUZo1CWY0nW1jxSjmwjD5JKsVcFKJp49f+HP5V45KfaFNXa7o7CSJ
NNnMePCsO+Qm7lWLJQvhr0BAZmcBbLrbhEhwZ0ORCxfbmdlZyVN1gPV06otf/IA3cB4zyws1gOkA
tnzFuVcWfQLYORT9TYgkekNdPLzjK2ndfWt+BTqxvWBmTh4wTvgqoAY9X8LTzRHufC2thrkmpdO0
8wmMr0MaczkHKQgPrC9L6piimJBpgVwXsQ/Rk5JYZRhe6OyY4UsihpBIb3DG/UbGl2KXFMB9TTgK
6K7poBMEhnBV9eonJ5723z4/Y/7Cn3KlLzxGdlPQzzxGJMoTg40Oxg33ZcyQOTyi4cZj+DxMb9Sp
WJf7cUl7LlE3q9dxrljrRbKXL5RI164TxPqwMC4tptsyXqcBCkklgZv9YUqoK89OczmkRVpty+LD
rqR1Fdch/1ojvF0TWw+ogEDWsDY0vLMqcA7bcEOe9Ksoq7P+x66mjAgFpqSW/y+p8XB0C61OvgY6
8Ut0EENYnas0nOzD2C35jo39iHNDNna3zCuz9FGtySH2CKLnz7SCjH802inhevU/Koaa2cOU8h2k
5IQicorzMlBVtUwH1Q0NqRIa8kAS58J8S/YgxVmp/fb2QzmVLZWq5ae17gIVcu4g8i7uEJoMjxB4
bzg43Atf+pKUUYKQ3XFO+xnNk/wddLGHgcZQwKHxkvtb4EY9jehabEOSsBfiVNZxHd7Yi44X7MK7
yu2Wr/WDO1zPZVu8v82w1loCuibR4pY2DSFNGd7R0Kb8RlrbQ+OqrrHy5mVSgUQ65eC0l7ar/BwM
wtCVhTOEQBqwJGoYG+fLNsT/eyP/fUHbEaeR33YzrrqLklzps7ZN4MZ4SkdPnA3lx0uAxGoCqpsN
j51mBS+jMQDlqUgtwU1Oersj1aUv1xnIM7D8y9M4cq+9+lk5ibl9AbUzF8ivl8j9QKEGWXh7gYZW
t8kctcQx7I2rGAl3FSxZ06efl3eTU46wk92g6IYf7tdTC0skn0DmaWMcCA+MoWZuac5Y8mxwH6NX
CPNKIOw2FSZ642fhj+mVfRArvOkKN92FP22YO+iI5AwTjVhSpqc6TRZ2yXH2xCmrh64sDodyDnLr
ZBV+6nCkN1tOMC5ngZCYAFLDIgGqutzwgoLLQfyoigZqjMqotL/DzGXdXogvrVpLaOJ0CFEGy3Rk
/1h7O2YX8DeQ/g0WKNeSB2g66vLp4H7Ie4BCNv23u/qsYUouRro9O7H0+SqzkzWxxFNzCvhPetEA
kdxU+igBfL6wuupGnyzvhh0/TKQSSkxdRymo9i51fWERTrTZr+uBMTV1jaW3JoajfJk5i9AlEpen
U2jcUZrnFEhRhprJWUUgOE+sfA8Solam/wHqxh2AwmkhAsDlvXci5eXfKCiHch3MuJevuMsxyl00
QOKMw2WGts9J3/D72TRSaGV8DFX+dZYrQnWjlH3sdyjy3V49CoTPzcTsr+is8YMbDnez32UuBISF
doZG3rM/nz454kgsqpQqp0zd2u409qMc6Gnl6IOe38UNar1KnDZ+Ud4BUpaSkbPtmrCaotbd9Ggg
M2qo/1apg2+f8k4kV7O/t0hVgkbVZKyg3fm1FxA5DbJDZZqjmnKVN8IiFMvHJI/P5Lq7tjmqUhNf
lVrxV9rfJ73gCYDB+URejqybbJK0U+SonhoMlKDQIChVbGaR6GvfAJ4jOCcFBJ+Or7oLwSAfDs85
U0+40n72aawKdQk1SrfSslfGF2CbONa1JxaBrUfL3QOr3xwifwZ6fY2kYDYYgUPl+6FdX8OQroWw
IAOGPq6xdD2a/dHRe6LKG4dR3JkyPt2n5ufMPlLjTFsZef45q/ALi43/J1BVJnxiPJio82EG4xH+
vFsT+wPyw0Ou3KPQs5sJ0lTOBph+H9xgyBWKOkNGrYlegKS1w1EG3DRb9+/DcsqJkGBhIwo2Hgj/
mbmuNT/oNcTCyPQDjhPDPDxo49jS/bkheygs1UZ+JduezhQNvUY/1Uu2AT3LMOLiqAser4Q8SQwG
eOHpriLNWT5GVFSQyZkkUDRa16/qIwURg23vaK+EntWNsNKAkJdmIjJqME89TZFY5vf2hSuqU6gU
vukWwrKAOlQFglIECB11/LSudlU9ao9jbgcy/SUFTwy6WV2wTpsKtImLbnTkWhW0Z/cpfOgYaNjc
79s8ndb4Wh/9Ij+31vgiPfQ/CeAYRHN8DPH1LcPScYwzkzScz1JXvodevoEAEfJfHarGW5gW8twv
pA8EAktR2/6VzuBZ4FiX/4/1bGz9n/ZzOMLI1InO9qBJfTfuCZlYXxCXRlzVWwDhls5gLUs1bdqM
vRicO8Z6Wa7ucnkJWV076eFz3DYsCYOcmC3yEjIhaAEqSzPVO2bjPKi/ARLkW3JbAHboj1a/xYow
/Sx5/0rwPHK0hUV4JFEEEE38B9tDcoHeX+PFfNViKVd6E3saehKK8hEbQz/4LxX/hF8KDzaQA5bZ
VohXnfi9Fhc7AwMetEQ4o+RFEQosy19zg6B+n72qwq4w4N2JXg8wyAQdE1xyHuSeY/z6ARnXYogw
KoQjT2KF710M1MsfN8bpIxlw40+P4N+1mM3xHabPQ29TjYYGVSUa20BMU4Y/EBrKbbbw7+wFni6w
50kws9GgMtYrQdulqNO90FR8Hj3em0idWy4gIY9auh633trxUtcYE6riQrpJQPqy/L7Mt+eXB2Bd
8elTe+vdKdGXFSu3pk8Onh0U8kNpLFteC1mhn/7M96s+p8D8SdVDHywVVp7MLS/alu3OOGeZ/ppG
7WFcqqEuzfUZEx4wxnvWFFdeeZOOyvKVIi9N13m2ZkW+cBLvqYbIEblt6lmKuA80T+T4GGA3Uthl
A83me7hU1d8IJjRlqFeK08qACgg7sHBMRU+MOBRqYdi3NpaDgotWg51wCmLmz2utPG6sB1eW9GrC
IPkxpCQrSw3CxOFu6xKWKZwNblpheS3Kx54C86yiSJcRRnkbewrGk+1S/6T9CPfVMsk6Hqg+A9SS
mEMU121vRaTIHr+cu4z7nRWKRSwgOedZgokYBObh5oj7HuWi3Km2XSJZY17OWD/8XvMCRb0HFG4+
Jk/moTrjKztJTw18svBcGCnynbYeYhBIqPRcc2LmdPkWnKwJHZlOVCnbO48xh2r9iicL0eaREw/1
bdjvN48ThqDpuWQYyd4HkJ8DOq/XRqxJ78Uw3TjWilssAxMIlNeV2z5LPa+I+MyUW9ljUr6n5VMt
nMIhrE9f3g6QdqBenHGDd49ytwe2aOZXWpeJSdxTxY07LvgiaO0n0gff9oO22zi6q0PDLvM6qdEm
Q1aMmEu1Fs3Omll6bRCmqYvJ5LAv03QD+kf9CgUl4VMozpYojBuie4Pl6R86CvjDV/fFPw7w7Kg7
iH7wymOvAuXlL369XKGNeFFf7l+WrDY8TkeQngok011h1Z8VIx/W6EGKpv8yKjRkTubRUtfC4tVj
JE5ffdko1lO715QU65OMoMu+rMMc5b1lUTfAzORjiYmNGu1PObLMykSFugU7PKNy3a6rqtqFQkIi
O2uFUf18h97IC1GmcJ8ZVIvhkqg2c7S6jE6bILxm6MbdadW5yY+2fe1scyX+w4Hi3G+DLdK91bDm
wbIHYLZopvxBTqdmz9kntitnZqNxtHRLHfU3GBTKiXx/xUADbJh8BOCPNElFOahgYUFpZ2eoXlfr
xEicDC11j+XFVM970FUTQlSzdphPWirF3nUh1ayxgBQ9HPO2osP5JIJytixdNBBu/b5FTI4V4vyb
+oKvz7agHxRmkBgXZiZ6rPXYL0lfaqjCqbum1tLoOWntGiPHJ5pHpNYwnPAOzpg2j4ew9dETG/1t
jiPfwvDB5Wi3LMzGujoEHSrHqS3TfkshKWUX2sN08ZLZfVazcq0ohVBrE7rzHseNPQnSLqzRtrrl
q53ls01DIPr1l8jnIkeB7kfiZ+rLiSY1Nug5iL+8o9Vf9aPEnvorj8uYB4rFgaXZ1nPranuhY8K0
3Jeet8WpAa0zxFikBgX5vsnK343N2MZL9dgpxobj16HeRmcQNW4OlTe+bx67Fzmvf9mZphk8M8/g
kHlsu3Zt01jqIQkDYQAsg3TVesv9v9ILcio4JI3jyRw2aszJ2aNDHe0ioT2WVyRUpKIVgWHH/XLI
1UVddYHkGnnKpI2VU7U/7AqES+Gwk+Q7aNabRSoYoO4QNZVe3zDMMhCRUAv8dvdvA+EjEfKsPt5F
CsGVQKDvODuyct8fRleKxK+smlVBtwGP/ftLVEhs8KYmn1SbzM+SpNddYHnq6oLpj4EjtbCfU1Fh
tGXOysAq31B3x/vvzL6NSi/M/wq/Gj8D/KwEBmBRUHCxZYVilM2fsMrydqggQtheLdS6xP/7jn3n
z5EcebBgmPwjruOL5J798qwF/IY1XY8YeaeHIoXtVg7TrU4u/Yjv6YIhbx3EBgMtxufoSOUy06jJ
HtiDgO7j/8IWmf2gDuN/nh4jfSg29GA7km1TvDhJ9vh1g8P9cCAWo8oE7VmxVlk0hd6VQjc6AaxP
3zJusRIE3Zbu7m+Ggh51yEKRNuxANagKZok4lxlpdJqU6msM2XjaPwHccmzZOI8tacPLLDrIzDNO
fnT/xs5NgmjJiVZsPP131TRFY3mgZZasHhUHAOlz6Q1pPH9tfDacvmW3E58WDBRv17u6cgYKj/pr
F4yNGcTjIyhQmb+XVJauJ2R7fIVdWYjz+AhrrxXUZJBxPFFwCwknnOm8JQL4F89baVOFQrnL28kA
CBMZmxt5GK7p3X9D4PbGZKr/CVEQ3cw725LqlXZ0bUDsDd69+V2rAV0yFUhN4A1C1imlX2Sd5Urz
hDwWMkSKwRjh0O/oF2fi1LM+12W6BTakxo0NsthvIpYiUrF0W9q1GBt56TM3c0EJSNFkmojD4LxF
h70AbvcxHKAmBbGC6Pt6mhhQX8cUQvzYdy4JYKypAyTxWZ5FyXpPSDcELXVUjCDWKoBRhDnwUKfx
7ENC8TUiGNf4GWmspkJH9A4cnvOxhEP92IN+kdNP5SoLjbSNkLnj2iaO+1+cC6aD3FGVOwEc1JxW
435CZUL2+z/kVjULo5PuhyzZrRibdFHwlTXZJAAEWiRPiEFrHmUfVcLKrxkiZMh/qvxmzqNrlyJb
ln59NOuv1+EJbn3fYzXQ5zQmNdOvFQt21v8MUMMsvlc8yhRFjXMcYdbJHMmSMaaOAy2r1E2yt90r
fxIOj4ZmDp8X60tN3Z6/6WPiB4WPqIWb/OalQ8nhj1bYLLoCaVGQ7PgZDEevPZVxQRugLWsUsXDg
SbEGmC8VMl6yfI+f2++zfOwFaKX07sSENE7a4sPqamvy+tI2pke8ubwZ1NAaFCeHPWKzoGspp5K9
+MLq1w44GxPXLe0fWr9c5JNwV9G9u+IvERuGmz1u4TRhANP40UeHSyBFtOQ7+glGe6e6NQsX89bB
9rfVZshstU3eCxa4dLWHLO6dJcA3YvAA7Tv2SE2douu4/2vyWJ2iqQs/Svs2PxMDpn6UG853hoBR
5EScAsl+C3V1U/SM6kJu2AnKZpH27gzewgQXI1CwiynjIO+Ec2fDTWpTl2xsWimKfZy5m0ckXeDj
cufsnA05FoJBGh2pDfdPVy2pScgDO/CUGz/xR9hBSvaHUnuhuu23525nosUsVs0Ah691d8fUugR7
dM6wlbohosRl5IRTjXQJP/oFQHcyDxKkPe7RRhni5HV8WQ2DQQaT/8i2aUPvdY7aLMaFhkWvW+Ro
QxBMCU5au3pbKskkQCPiJkWUgxjr27gFEVCWXgbYPjwo7SiPsUE8sVbAHzGULkl/eObGhawM9/b1
uDWCwcVHV5DS/+itQnMhYAMPC7dzkPHEPvxGvpdtfv1Y1MjdKJAkygMrZqvrBKZuviI7wNszIAxH
verQJDGCrp1TBnx1AKqL/hY2RL0Jwy6jeewWrNMBHfxIdmk5qrzgHmuq3/1rUrmiqfz1l9HpiVFE
HWaRHLanM5/X+LvBMNWbPS3NFBGy/uYcjRETeaUC8WwDUnssM03gqVd2SrIlbrCy5+8mYpLZhhLw
DKFWNV0tSbVyGvB+IBYNaS9YDiZtDBQuEkNxpx6umFVIiySGOlIOiAF0GdHB9rnwCYMfdK0gdUfZ
GpnPEsWlEmqojhaqwba0AWqOqq1xgTAA5ubF3NHJ4/mI++wbzaE+piFyplfDkB0b+o1/gnbUpol0
zpitbSc+cVyU0/EDjohEi4KYWQUNOQppv/M0ZyY4hway/NDjaWNLNK9plXJ9RSRscDNqOaACDU2r
oJ0NEgJwRGkE8FHx5oAn1rhKv4sd0A9WRJ5D/KzI+LCr8iJY2mtAq4h1HAy2Th0UjTdA07NYxJ/9
62WYvSTeV5bph/KPc5UYRmoG2eDgCfiyTpMSk2fOmH+XG6b/BxTwwir3i91KE+ZRgn9pedCwcgxU
d9LyrdChlJ8iAOS1OaF4F7pl8tgt7N6UCCkj2iNGA9C58/1RTGqccBbMHfiHY0bVj23P7wmRLnSE
Gks3GOXcLanJlpE0GycStw2+25C1nPONUAgK43LXaneHuEWsGkJeaVXK3VP6dQElGMPpCzjWrBln
8Kr/raAsURgYkATQiyPjBVyMf8XwH27vhk3z1jypJK//xySjuR7LBVOUOXQogF25ipENJKuj2uXz
1HaWVxhljY2TmnrqRWcdgaoje8U7MR+6cAkNY7dBRuUA/PX1N9+s3zXXnOFzdQb4kCM1e4bBbHBU
8KuCqi0p5884iBNK2LagRKCo/fBlZOJHQioE4ptmzfmfO690u7dsOO8HEXDlOJ89JrFwYvBjYJFP
eSqVJ2aPJOSSZeFI1+tC0wyOxNb9Le45OHKanoWhGjqMdRi2Kciz3rAH9faT+eeyRzU0rd+//9ou
XFqSoCgd18aCyzL+yFxTlcaNfeFUgGePSlrasNjpb2MLGdQYdH3vuxHOVZsni829ebBI3xysAMac
nvRp//0za51hP3hJHAQfOzFVCBqbkX++D7xeXMJd52h+mS+iGe++n0dGQ0uA1CnWpGWSm4KThIMY
9bavw4ze6xJ8dvOTYoihQ99huFJlQnyX4PX/oNSvJNrFH/QtNI/RFuoPEbwMokOFbrr/zl5YIoa0
RQ2xwQQ6M8JhYHnmSxeBifTOt5RUyX5E5mDSL+utBk8IBb99NWkouAO26xm0meahmVTqzD35s8Qo
GjE5oMB8ZZZDlmuMp7gxI1bXvrrLoP3ilKXWRedCEps2O+WJnlTiFW2iV4u6au+eEfzQdsZA8zCx
aAn7vERcnipAy8GP/tLPSoA7H0MQak0F+wLh3q454tzqZ2je19HkNzEhKNu5i30LWZ4IKKOU1uqs
JjhH8vzLc1wvcXBgAkJQ6IP2xVaXEZ9vK6GWiOoKcUu008HmkB9CJxCPaI5ZGcLQUUlz9zisMer3
5v0H53iWzBuW2RMR3vzmrRNvISTqUf8lZWOJNSuBQm408gXlf0smTSa6raa4uTRR06boGQrC6RqY
f4TlOIedR/FVmCiJ9745WRSrKDD3tGl6P1zg0vgdY54t9qSHu0SXiJqhTY5luD9xxBLPgtqbWnQi
UKbXmvAUNCPrQEjbeybar7HgM0i54ZQv5Z6IKPeZb6dYEYAUjKLrQHl3b4GjjbN8WsSjKq9Lw34Q
OB64W6faQowCVdKdRFFOrFmUO6SMF+OpTw0vp98amPSf1zHLVbOavJfN7GRvdBKHVI5PfLHSjGrg
6rSvu9VfwTwkWXjRRg6UmmjRjQgFYHn4yz0Qod9iOagY8VijyEubTV3BxfvPsn3IuJqgBXOxj/dE
d2aJ7y+YAynWcOwDvOy8BhfRxbYDqLsmQJElQSQiH3k348ljVTSg4DnrBuKMOStdDDtJ/NDSU11Z
d0QyTyIwLA69uRZRRW8rionizjZgd4VLmy7SFA/tHFoX8wBGAWuaNeqn3kDr4uNaInkTJstzo6hn
vaGp5YzRhvbJyAF9IMCZgvcy8F2MPWwal5lM1i3nP3TmQUSsvkBLhtlAU/FgMIqiF7WRbeoAA5oH
EmnHK/Ck/C1MnQ/6G0a/xMLQCCMacgX8pxoWqMl8BFZIjnlz08ZBxUheVodZncP06DUdS/2EhpNn
WWrEgExBHazwlIgjf485hdAYeR49DpExx6DVKynRfqrOSKmkpQb8b1XFmnc+0ygnfjtxaMDtm9ZX
XMwB/xL2jSveuVmGzbNG4KEDUb7rWC1634gKQCskB+nijcN45zcAGoDABc4m/J4d4bC0N1VCxyZM
sLrV7YSMuaZyapxpbW/pzFMq1HgOrRUro58IrCgMNVzoKFneYkcvaMKmLiMpwfPE8loKNvdZB5Xv
RR7xTaf2rcztaCJ5Nr7XOre06G+pbXDX+zYHJv5+mrbts8tpJMpoEOA2evmMTQ8/3se9tpgjPe5x
cOgatk59KKuFEo9NE0VLc/kc3NvUgL8T4zVlGGqq+rZnFUIRAgBM0RcIYYePHt24DKxnBFVNrYe6
t1l+cdMYTwFtrQ94Qlx6+I8+LJa3CBRtkU+6CNNey7uT5e2WE9YRdA1N1r7HcITx9ED8onNzQfDt
G73y7r4jT65RGoHhdDGbYF2eLzEqAG+Xp2umIRZCXDMSqrVBgVH79f+9M0KifGwj43UI06rqs3CI
YZyRx9TPqkRjU2umKIc7fCKTKIAqeYnwJmbG3W7CLZfcEDCdZ6f6zqrI/EEbshmc6ZpIY6xOBMcp
sSCIv1UfIMbDX9XaCAklqcHeGSWsv+z+s9APz66xeYv1MHrJZtmclDLwb48YL+fEDDdYS9LLROcL
pTIdGWDdein95XZtv8FpMl/1fAVeuUJliMtDn/O82EgT/F3OPiqtLPx14sU9Ef8qwfR1mO6Jgh4b
7GeedYCLixmAt6hm1T9I738h7/ZlUuScB84SafMP6buckNs++oPehFyvpsao8fIQ4TkTt1byyvqs
93cgr0SnB+NxWmCIi01RFaT0AWteO4Ieedl24Wuu952VvuxnvdOLvTp1tdj1gZ4CEpbEaH2+e7Db
T1X0+v07vjGbSZQjR09XOfAsWr22Wq4lolDxOCyUc2nfcQOM6K0FPKOL7UQ7qnfWTKpmgI1GUtRy
L4TV/dAUsWILQMyMxbG4yOZ8is7XJnpzwP1wmyB+vqrBX6MO9pEKTzOWU/SqALhYdyJVlZJg6zlq
99eKr3iYK+jVNOreccccrCH8H9Tf/tXdLL7CqLZZGTjczPKGLpShaUh5Bi//cqy/pjYop9ZV51h3
WZoL8FZ30QIu1xlG/it48XT0y7OAEaCINn4hA1GcVdG334MUg7o/Bk8reZ4G5nBRCFxrO7DhpL2r
cBl/uP0LGyTKW1HebK4ffwBRM793eGoe674uUD6PvIGCAOeEKe4IvoU2EYuGKuQVIx2y1MEKHGf7
DxOM/tJmlPlaDCVbklpgJgFvBx7Rm2ftuh6Y4KRCnNsQNzgRFhjrPt8SMbHWZmBqjkNb3LWLDaqw
AKq5RF31+muOA6Vid9jTQ8ZuJPEMvUKur21Kt+5Kfgpj1fGGqcorM+Zs+iWXRAl/QZ4v0iYkISnZ
4A0Xstw+RnQqgcNaFIg6w06tdCgXk8CgU7Q+BFXLDBoEhwCrT7rQM42FNZ2PMVbvVhsdlKSSePgM
2uRjUMNn+C+tJXf68fqtgKYIypEfbvsNfmeb0IG6uFEUFWYwonknO44ADJ979mecS7KSKaplocSH
ZtbW1UHhU1PdkCaFa45J4K3P8cpsWF94gAMfFyKO8ADtnFXI7ER2+1AYusQkC/E85jVeh/IaiKCH
fSgTlNoUlmyNj6tL5+sF0288SfiKqQtUSHoq7AmcAX8P4WIzxeDl2tQh3VGJrqn5S2s8CVjzAN33
BKI5O1g+341gUb3bo6KYY7E38LIjbf+k+mAQucqgxLRZ222eEGu9miSnIeNQtn0kBwaxR2zu0IaC
BOFac5PYbjt4UF4ePLpECh+aRouNdMqzsOnQttDEzSA3KnKv0DJPXIhVU53rcJUDNXxFV7kkCJgw
ssDCHLOgO44RA2r2acWEhcl3mz/3N+aw1FmYp0yAlwMK0YbT7i+D3a2tpzuWVegdA1lSyv7+5Y1s
sO4ueZsXRw+B/mVmAicQGwkgSv+LtKSv80W2VsOL2z7DzylipY3c8GpoOUZIKjFv/8SWKgCCeWbf
9wRKdxEt8nBWh27xGwEEbwD0iL//a5cAB16W0Fd91k/cC9R2eWy2tIPllQr9QR6gQ8WaKlUkzEIc
3IZfbqBeUit9yvoBJpKAv3/WTxqHTF7u466FsGi/ZacuYXo3d4OEHR8q7XD+62iihjC6MfioDL4O
wdzJtRAl8VDrR84pOtoRPZQbtEvvpENBv6/+d5t6RxW2GIfau0+QheErYwKvD4nlbSDMeeEUWA5N
/Vt7pjg+lCDG/khRzYntfqShajJCu5sOJQCbpZdkgCqbDPG5JzcgfJbHoMMatFt+xQ4V7lZmF5gy
ynq4sNiW7UyJ2EQ8yOfWdvKp2IIm0kNBYoqWF4C3+Z6+RiWkddkmq7HLrpiGKjPSS9ikjBTKL6Zr
bdLO9zPyqrqKnK2sDRtBAZuwy4xQxirfbb9/QEp5a7keEJnRw5V47OgdUOZx0/4VfCKBvV3DQNQp
+qCIhfbqlYN9PLc6GyYCzHdy2qM7b8eAV2jwSLCOG57cc2ycvhulYVH+BD19TLG9AoXrve6Rkynb
OYjirF702jbACtF31lQZUQ579ZMKt04/ZCGuf+Z8wGx7/Ke0vtROuFEC9fjuh8dDYaA/z/ISXQaD
33Y3p9xhfMI+9mbabv5RIbnpiMJPtz5eRij4S6M+TwD0UvHqnP2dQAp/SoRmhXVyI63QCwS+6Fsq
iZ/SLO54NXEZwZs1U0GSNQi+PCrqWV5Qyf/0+Qysg/JZMuo2n4AIsDWuN6t2LW8S89haAKgvU/St
s2+dBuslnmvB+++Sl7SuKqd3HpHqa1oQDtnLHbwqBbs3kMWIyoW4cyIRV5NMCYyH/GchvLyg6n5r
jFPHVbPB7/6QvjSLPF73v0uHK+hUutJ1VPytiWK0b3TMY5sQJqshc1d/9sfoAtvKvHPLs3kO1sH+
1roI5vS1R1wfa/G2DW3Kf/e9QKPX/9QtapqIL/tGdGNgE9B5LIIT2cXdRZ3ceKiWSsKNkpXSnzLV
5IaPIjLtEAlNsp8W6Wj5K9aBnBpFDLkJqWrjClqR/MEVfEVRIlCe9gUmJYzCnZgJW4Ponuw3pKjz
uLw4Q4j5QSwBEG4nzEIgJVbB/HqGDwhZI4emcwKh75ySYy+zs8THVsCGF+2a0z316P+OWHtbGRdX
PTSN9PA9tVSawqXlBlLq3UbNwLYOmUhL2l02rVj1+rh3gXpYYUnkHcD+OnuGHtLeAt3PxoIOxnPl
eQnycBjBtzdqNEdzzKq4mhMOyxEMdetn0ky96ei+EQj4ZUjmtiDjWpYplUTHRDVu0CQGAKtTr8Cz
LjxMXT82jN8HsR1O0UceB09YoEeNovUIkd3nZ2x7furq25gYuNyB9346dNmCPOB6N7ir+koeDIor
/zTtYDRJh/Hqa30dhNeLh5iAKuPllZ0Txj9X4l5nC1nxQ9xOkP863fETSNm2xEXmcJmGHnQ/ANL3
rdJ1yGoSHyBusTMiTosnLaMo85avHL42xdSMt6qKdb1Z2/u50OqL07WL8dF3sSFCKHb2iQ6YVeYY
aDMC/colDxmsdINT1NKWQ+/Vm/7eaKRfg0HSyahpNctfFZ87SOwrRvzf1hddMZaIDbiYIUEHIhDG
KtnDgC8Fu65TYypNBdRW1tl5LkVxm08F30a5pi0UnG/pikkGmQu/u1O9iF/vnRaq9RoYnVIm28AY
+XS5Y9J21BtN/KCgCauY2Oie55v+KeOCz7iAk0dh0xanLTnF19CKLQftKtyqZu580GzDtkOsoICk
s2ff8l4/JmIbEf4tPKfJVxZPuMRKm60fliXj5xTb3pr94NODlCYgL8LUSkf4IOonw7UnLOjI9QVF
8cf/k7WYenyP3Vc9L4OCKeTVUhsjPkJcZ7BQn1hCpOPaBwUqiFj/eoPGPn3ep/hoH1xWeU6zpOON
8c34wl2F39wqH3nzJ0qY891u27WN+Mx79/2Nb4w4vTkC6ZHQ3ooF8Dm4FtFdt+hNOPgIbRZ8Sabw
ZFgCH+rzBBR1EIcDpXQc7hDippFmamGBUtab9hFcZYM3ycRfki5TiE+4kEVcfpH2a8v4AgViMuH6
fF8FSXGKC9Q8/HCBFMzJpotQQRLOmpXvQaHTcZG/Qth6vbhH3X10F99tldzlSQN7MH2P0U3CQ94z
uSoAR0E7Ol727SUSC40XnHi7PAbOT+bBlIhfKKVlt870swaIyz5eLhgzcq8rUCgVg8DPm3yRHhgz
WtQrp/3ruG4CIFGasrvIlmPaw8Ms3562nh6oS/h1HmveCWMT/gi9+gMTYnHCJTHTfhW8wB0EsNtb
45xWY4ruj3udkElFGhcnnRqwPbzfeS08l3g6HHoRPXenPlmCL63rL3N6ksfNtNKYlWwCL+3p19AS
FNWmEeJeJ0rgs7o2lMWy2HU++R6EuSvEtLCZzqT7AQCUUnhV0PuoxsRoBjMVY4PE8AbR88wmWFbv
f6xNuIofUqgkERIf/XoFANUPzeU4JA1e6VDIe6R7c5G/32LBuylyKaKkLL9M5yC9QidmiANqKzjS
fvkddLAJ/pwQiPk1N34lWDGqhNCa0lxRJGpWtbHIlGI9eBAsQ6FUJA1q5PvaAJFDMjJdLRpx7tU4
oOgNlxKGC7v0kFTHCoVwn3hQT69aFqvSnLNDDmEF8ExXwWDT1uVtVfdTUycNQZanCARfF23WN3zD
H8QiBLUr4gN7H59wMXn2IePP/5czxNce4OAJ35nBHRrQ9UvNu0BGGT4eFD8+FAt4+l4qxs2WZYl/
rNGX8XleMQbMmmw3PVhkJDRPHnVD69d8FwJHwYWY/VokK1S+X2+MUdWXHW1QI/HE+qIGhaiNmL47
qH5E6E4YDgesEzmkf9pi5NDKxNkiJfVTxEimSg0Pfy5r6EjZELTco8noS9RgqhXjNBReMnFKrFvZ
PhZaNCGsiw15I2VVric85r7+vOjWLrkv9H9+Q5UVSD8PobUB5tGQ/JRDwEgxyS0xCOqtAduLX7bf
aSwm2ER9RdAnt+mOhMfI61mbmHG+b9s/lAjgVWLiG/t57SYQnJImUl0Y9K+tvBq0r774pUXOEy59
4CSUBNxBWuHbwE6/nmTdmGlO6KrS6l7HqjQSrFlBA9On+0l0wvOEGTZsQqVFLEBE2nEG1z9HasmS
u7UZ9K1ZrLizqPIS/Ueoai3uQYRTDRZFzBcYpdIYi0VFtppFozjg79SrGUiOvZIcr4cLJ59DMB39
yz6xFYoUyrx4u0rx325vSOxPHm63EXOVEPWpO8c2ZXab5migZEayF9PVyUqHmrgKwDJsuJ80GZDy
CQM10adP5ySmvYImsiTo23fP+UOwvoNhDeRan0f2tfEnmbFtIbnuRYa6rURVop1+dRAKaMDiWH7A
I//4r/o9F3NQYtQ2kZC475CfFpslenrK+i7oRlkurEoMhTMkuaPQ8j3+tKCnKbHutrWkvTy//Frk
DM5nwMeUXDzv7YBSFTZMHswgQBGcxpoViaCDuMlDFXJ2+SxzIupo5VhMZ50vkBacKg2s+lKt6sba
16p/qa+b6xMfr5mFmml5l+CH8C2XKJj0KKPhucXYHLPqifD+2E95ARomzRBMAEAfXVZ93hGYkdvK
xoPVjhLV23jNSTNASPTb59UYr7XthOh+CQliob/BZ7oGzRoxgI7d8ImOV/Xv3JLlxHCtk/LPu4NP
JqLooWYMblKlXrTt95kSy85M+rcQqYLpn2s++0S/OzmnPyqKAiAsKneZo362RMxpztkmOWKRP/86
Fy31Fxa0sVY5CcDnE/xHq4mK14bsryVnKaQ9rjrnvBkSCvnUDwbVd/P/kBtRwedRmKwL7r3oeYye
KDEySEjg3X6FFSiFdkWwCFDtc5pT/ZOfCtAAmJwPKmLDgJWkMQnaQ/QCyBPY0299TZBDZOXdA+SP
IHHDgOy9XbZPNqQ+Lp4DI01o5w7qhvYjryeq7LQirwrsxrIJO2oMjeIYNjXRwwJ+zVYGBdS9aZ2Y
lTW59ycGZLQdJTQx/H4EwiSsnj5cCp1uRqU2fsV9CdWcevxKQhdXYOkJ7IUnsgxfZXliGHtTvLMv
k9hbcvLk7B0ojSFrbXDGVpkA+Zae58fXwdqLBWIRc98rAFWGsx+he2KByF9mq5vpnFnOx3B0Ehmy
RaxQN/o7tDMG+fNy/OaUYRZ3PkWtrx3q8UMk/cufbQmkQ/hpQWKdzF/TMA6CH+PnmBiGKA2NwYsN
zDaZMI/h0gHQuCMC0K4ApFKy/h+58P2DGbXZxUv4tuyWA8nMo/3rAWkjnr9KtjsRnwTmd4e2ceH7
qrJoe0hyJ9Fee1UlSwRwkhzl6i394eZxxLVOLuve0bv9s8cyeIVBh9VrJHvoOt5vwgTpAkBoRqUU
9T2f2TL/4HD4tx1uC1mx50PlSv2FIdre6Nf/9KbXoxw49i2XC5ncWtKnv41KUOZ9KclyZ7zc+3cY
1VqusIlRmG+Mn0KBjsgjZ9i834nAPgQpsXHfIbyc28uqzAtTHWmHN/JfiVG4KqzBAlMa5DKTBlXE
9lFBsNLKbS5PgL6FQwqLoZPsMv1chYdNPju2SJLcDpkEy4jaxcwuP88sS31S17doZ69vDJhLhwaU
fEGe2w8KkoLVRR6e+1OOtz4TaI1cg3CnYXQgBwRdIAQwG1m9ckOBc6QPaK3IV6S3/mh6GEVtOGf4
MPRhc62EEQy68PldUd9LrjGPwdoqP/nJmZoq6Iid4pVj/9srO+pZcnPjW4sk4pfRII485jTvE4yH
0pk36GLVoWUPTcgKNPvjDV66X5d8BhgjLBzCyL4t5Y938IHyB759+4Zz5ETeD07o+ioXSVc8MEd6
sdoWHL1SUKKhYI/HAjjP9xj+z63pRanioNp0Yi+EmNLhPzGfZXXys4bGJE6WLWCgmw4WeM4lhGVZ
np6TzkB6ltD72LPyPBn0EuqInAt3O9I4l11c4GOsMHe8VEfloS1+07ff1SQs68jvbxdF6rgmwy18
GTPT0Wtj1kNfpJuI1cjNoLY8SzCjM2Rz2CMjJ6IjyyT1ErWsK8e9lHH77OZssmUkQnkekCpHDLr3
wObv+nRLuYmEf0UsyCAOc6pYbhoOZNIk1m1VY0PwTcZaSpNsxH3fqS+4wex9WjV5jlJ6hTG2hd+0
eNFH6VDI3HVT2WthJzEvmHiXaCKM8FO6tff4vh/mlBT6rRQZa5+01eJ3K4m35k5qtv7fw0Yg0YbC
GZMXLVg9qZirkK1hTlcu+kyrEXikfogUqqxsfUnu7YKPxcosAPnM1fxyxiGMctw/wdEGSYsOJNr6
iN6qSas/M4OxHF4+xc2VzJoTjqv8lc3lImfHNXCWS3zpFjaBVegwfAnr0AlLq8EzSJlEfVEjtNZW
K6jM/6MJTPgwt2RAD8b9bIM4jNq7GhOhva9FND9CJbl/TZuKg7z7Qnkpv7lckoefRcbvrusAmCu/
XYlUmpwZRo8CuuwwtfAgzbjF7Ut+Y0DnnBEUyLvE2Dd5mr8ndK7cSKAhXrkDdkHYb9cKr/+PzfVL
/aNsscSv3vfv1mlHJvDmx53B/EIESE+CvcOu2IMxixtOFeQP3KinBk7ys5PRtcV4IoJ5j7PGsmFK
V8cCrNM9rXM+mj3eBz883P0icwOVsEN0T2zOJqXaIXx1fpe6sdiU97IwaLw9cJuzsJ9d4UD/4Y6g
prwTYdeHxcCWQK0QNIdq07RnTnBHPn8MX2Nv18GO3aaYT0mIabSTF0qbhGWMiMZnUiKdjlnY47gX
OM70U5ZgArTjg9at5me9n8fxO08UxoCHBd3qXHVzdGfaT+Fx94Pf9oX718lua21cqfbDBK6UF4Wz
DxER1ZkBbybJ5itc7VzcSkbMMkRbfdYVJRWw8QlASzmfvBiwv7YKE7am+r6ud1WAiQ4NqSkSk6Mg
cYENX4rzoSGuzPjzZpQvUI3Um634OXMoZG4xhjgF5k+H21XHA5qu0rm8FfpenfAgPToElHIMSR1s
5nmk3TyVUpd7HSL4Von83VypABf8ziCoS59WSsDM2+185oE9ogDgZtxEZX4tRaqDimLDwwDT7HiH
P+aHwoQqm6IshiC2USQJ1Et+0UwVrvm3F8Ogy19jz5RN6wLVNn0DQwPxRBj6Iv7KJd/coBmMQQxl
ty5ujEPo8tFYZR/0wDT3TQibvtp0tvvN8L+cxiyZ1v90RjNevKwQxNNmSSuOQUb41KDhqu2a9Zxs
hmbsQqJg3KYVfcp3OZTRRdJcZyZKLGAe0xcOef/24EbmX5CafU5smIJLBamN24ziKWGB2O3WaJHP
BhkMVzsttvBwaR/3+mXud65BiHdvqVrG81K0Xvk/IQJxke4ob/+BNBj8Xk9q4rqN+UnptLRvWh0a
qEHnoqdtcmvw4ZKL3TREQDYGN3kzPdLhzvlHybkbaAArj+XoYDmaTWeZ3w+fe2hL6Uu02gpHxTO7
/r/FRkeFxwlnYF0mRxdG2Zbx9iQUNWE0zXcSle6UKibdWVskNaLLdxcuHkkxYsUTlARrvNHp1nsK
DTTwn6k1G6dzxUCrKqzZFLox2Iy3IlCg9e1Zhv1mpjaFwrXH6qEK/7vPUODcnJYCG0uYoMq/yNCz
KMXXaoo5s94Av5E4k1PFNm6IhOF/5AokQpQnEj2f8XDRFlCNj7iQonavkZl9K8299gECVRrvu1gK
1LW/2ZFtdYjxngVQMwTIpPWXT4HVNTQJ6nK0tikjc55Ae7EVff2WEZWyyuRUuxUHlse3H+gGYeJo
1oJ14sY4VRHbNDuhu0vwcXXctN7Yuy3Wij4r4KLScRk1CurW32cYP3aKP2+nQ6w2kqtKbykKrHd5
8RGerrATEWv+s31su3Z9XHDBeyrbBl0oOffpU+Zq12uRcFtWcZFQUgvB7MSgShjjvbKrTDN5QMVr
xarK/iu44CbNYJt32LHhYSJVWFnvF9bqSZd0pYF8ozknCV8yqS+2G0Qt/brC5lWUun37UqbcmLPa
CqkNwKcizXcyyoBxWiJEzutvxhBcjEA6Y/wCDvf6H1jLjbXszioMEbfW1PKuM0aRCnAylzGHvLhE
eM8VPQHs33R+cXScTsasjif9WXXLOGno1jn8lanGMRzq9P006yjs+gJXe50VVjyejfSgwPSVERej
PylGkoTQqG9BM2JGGiNQgU0L81CC2EhxKldjzw1LSnIJQRO8YspLXrUD/JWNlb6kkLNcZY6xHsMm
HCXK7InmJRN0cJ6GhOujMg9ZFbnFkcLGlly+/USY+TJ+xAJI2/yGUokphoWRV2JUiFBKxqQPPM3n
DV8XINhaSYVsk02EAmWusE57l/WwKf+FuG8qoOM++nN65igEe/v9Q/ZRYI/+7b7bH6tVE0oDqqzP
tnB5mVlp60b1w7IVyZ1kJk5V2hJXB7wuyWTMnfFVQiKuwDjrztw2gKh06DuImdBUbaZm1D+kzrul
QbdC2FbRN3MKIUtWI4Ah1T78X6+dyncktvfW8oVn0LbohznpTQCjIz2TZ/CYJEdrOK/di6EZM6zW
E5Xo673SovitoJblw4+nTbI32xu+6sKGzLw7YoTV1F0GE3TeTsfUKcEfqR3sYg+uKkIzKC9pFFKY
0SOi6Gc/wXd5jmNU6kXcgfOcsaHG+h5Ped+fF2ERTvVqutQO1c+/c/sXKPG+nwfM9CZZypzWllVp
+9NuQX2/bh9xlVy5fJOhOdEjzrsP2ZmhI039mQFWgB4Fdu2RvtVt98okvipPNovmGmI/N+XS0lgl
kbL/0bzWcn7O4DZbOA45bKfD17E42viM+Jl3qaaeWcqHbbzwPWCBCS/Dcpx4d4vu9O7nt5OEynDg
RTCTLanmtsXl9/48DctVawCRPxiRp8/qR6ZdelI7gKLXEWXQuPo+VNy17EzZfWv9Upuvw+pCpGFZ
xsbalwhpxH6sobq6uuW+5zJqTPzb+5lRIamEhrUmBvvgPLfzqmtWixsx3VshIC2xan9iqDJCf0PK
JDpUrBgorzOeAngkwO7zgduEnWMQIktDwluS3NX0wju5g4g4B7TyPPmlvC8CJ0YXenp6FN9JzYOX
ZeKJL2JXKiNqQ84biokA4q0JmL39Cq3xBsH7lURjkOcItTdoJ4YZzOwxcc/tCpFRXds6lDCR9t2C
946RFyUFEb0YZqJjrFRMYbA/MogiYd/BXsliV06nrFHpzgzRYtneSR1uBMP/lrmavS4LNSq0JSfx
IELM/i8t3N/fOg3EP7STHTSojX6jdRcNG8ppoGK+v7Dok3ec2QdqGaxMkyXoLdhLKGloTpK9bXP2
K9AurHndckLnC34dv8kyEfO7Phfc2ApsjvplPGwEVZXmo2djWjvaB+i9ETEn26kacerTkijNChXk
sAP2eIFW8JAyklqz+HLQSeqH5rYUuf6Ras5Ef4L7Y8DKT9fbIXipd1uH8BPX51uyPU8Cg0XV570j
DCB0FrSgCLmTlaLTPT06vxONVEOQ+40HRzK7W1PNEsxQqQMTpNXHBJ9WAIYmeyK51dZZK4wmlpSJ
HKdToQOSA70XzWkiinGlaULUedhW7PrFQeDeUkqYrDTQmBluhYBTQ1w4zH+6yDxK0Nb6+ib6lMxq
dMbPvvHkWGNZp71o5bkvL34AWgoPJTfdjExw1ueh3BhH0sUbvRPFzXSRGLiU1kivbaw1xgAsbNSU
4gYjNVcvocSo2oJQZCajjR9oQQmSAYi53TEiYfPQD7WqY831EBScs8LnUSUcVyqnQ2t9wX+KvaTF
MJSCmRNNLmW3DlWTLcHlpE+DmYvEkh2JyB4Xz7D8WEqyrp35+0ctz3gY1dlhjTMKNA7Cezwo7Bwj
mf/4Sh+DKWdS0Sjh35w91e7QoAJmEXR/1ff2Pslw5KTFeYFezkNU1tf6gsSiPPcP4v5VOK+Iv6er
xbGO4hiohl40lxUEP+iYLGF+JcCowfovcy7zGnb48jBR5natp5dSW1YxOhXOzsZ7JUo4YIRkFG8E
ZHCAdAn1tZCJxuORh/APFihljY20VZgqQzpjK2aQxuZhTOxPASxjz6YZ9+2m9fNdAk64Sk556ng+
r6FSYd7QAtjj5eH2JytsXmsEhzxQugg2bbSPA7FliXtYAZpTe6778XvkaDdpEjyXugBYcIUKaaUf
9Nq6ZK1mRbyvq7jUSbri5+Qf2kPEjCUjxs43CtPsbmHQy7TzVqtLxv/ABUtepKUMB/jRd03LwVCD
+iIuUyBdJ0vi+AgFjoImLm6G62LFhYxdKskuEeAeQxtBy8ZS5sKa4xN4UTBHX6ovmL69UAH0bvfX
a5A0cp5J5CptvYmB4swHmC4mMI5y9Go+5xDBECYwm/n0WmzCcCmXNLV9CwyuYcTBQhOPKIuQRqpO
0kKEFx3S6fZhMXe2eW6m3NgwuP+JEGfcAnkIM3HWMdHZ7AvNOZr3bHcYKjtUxCdpxfTbS/9Oslth
Ei0Jp+jIW5xHNNyJnr1gMo1JEsESE6O/9Rzrx9nxNZBQ+Nlp87wwMlOax2KiqIJD9yZ8oXtvwfMK
N4//nNJ4f9T7WN6jTu31k6PI+a+bcjHRdtB9xDfgOmX0hgJdB/kmyLBZbaFdYkuXQlnniw241JBK
tKL665rbEpS41C5k0N2x7Es0eo91+gTll075xIchMLLdzhipcRg2/EGi+XD8XYv5Z5PpMcjp2b+G
WRjtU6Tj4VemTdvkyc56e4kjtoZjubaFe4I7oB9Kw2AIc0GBIIWva3auQ84ecNt+Hha7X/bzTKDv
UxdrElLFazdR2UUabxDw8W+qxZY/cAw4sEmjR5L+YfGM366eXAw2MnawUpu6A19pL6B/IoDv6E+3
ASBekMcBwtK/TsBaWr/MmrpTeTl6CnpAKLiIaGqJ58IIAUUw15/pYAMvLopRh66fyOuHj9fT+shJ
6uBJ1xMFRX3MoiBJcaSHo59eiUO1eVxr7Cdyy1S/AxJ3erJDsecSrlX1olUDVR5cNVSiPWiH2hl3
9z66Bh0o3Z6cg4V/5GWwKbjna66PPankfMRiShABDES9DYbCAN/qsB1XeQofAnt15orY8F5UFzWK
evUkxoX59W7c9StOqoWdl41MA5IuanpfPwS7s6T92SuvYbg6h5loCxV0NUnylvJoHZ/DeeA4hEgY
uqc5hku92vQ9GIy4TfqivMFS3TqUUmM053yhKuVl++RdQB88mPcruxivsHZTDlxkf16dFwErOaCi
P+q1knnmvmBvFR7NMgI25bfkeejidwu9ZpX79cC7NO63VPySm+d7w4EPLVfC2wAvUsinsNZAYIco
5mrOUt9MX71laUFIvnz7aIw9xjlm1wJ/HK/zqvsijRDavDCHG9HuKcOXOigFMCgwWT46cn9rvU4b
+VxbUOs1xYr1UBlC3GYwpTr1/56CUzH89QX0iv+EkoDKA+Bon0NC9gLo5Wbmt/aa/vGoPkJ+r540
ovtVkSctE+hQDWiecGxZhqJyS8FMrdzOIgCkOsGbG85Ad/WN+IEoTuEH5KN+22pAzcPjKwPeLmwH
aLCFfNlM6PgPvIb4wg7uGeORuXLxh8sIs2mNceOfXIN1m5I6uaTdiEAYSdFwLbOLpacS5+ERFLgG
ncNwvWU266eUq1Mw80L5wiFYIGYhnd3O5/QIYnumkatfK9tGX8rPLhDxKZhgNMgjDktlE41qwZtY
M/h4v5+TGTP8K1O8sEnYvq8pjzpElhg76KElhzxp9thOtfn8qCjGnode0HKzjp95u0ftitZ+JLYN
OelZE8Sbzl/kgal0TPUV7CI7jmzB6zhgXdBIx3s7Ik0e90fRoTAOuHp19m6d4m4gkfh9y+dNCpeT
73YyW8isZP7f1FumRRJKZgoYavqO6kOrnoVxP/Est373uvFPig9ugnBEpsVky9u1T7NAoEDNB9o+
jUkHmIFjoBmt5h8GXJEWXCAqHwy4xs1D6pC0ojeWMKz6X3ATLKAyiDvMov6zE2Zsz1ejj92U0RXE
ZJ3WzEnla8I4KeOFTZTuo1cPGXn5Vd3pKfuJqQT397Iqpd4FKw/G1QOPX9MDIIRizXEhHBOHyJfL
5GLBKhBd3zmdwYmZookTg1u1/gJP/7xZs2eYGTpa3VViRj2lvQpjM6zDsvjLh57fpGZVYr2o/5T/
HryrfU2tr2RLKoXHh24ueP6TsgCYZfiMv7RzTbDaeuE05A79ujEd7qmXla8ecVgyRpu/2kbZTCCc
oOpDSDhokB45aIKFD1pXogrLynEhYGW9Iyb58PAH7lK/lwiCruqxNF5pgPvKd/QzBhwhwDnawE1Y
DVmaM3MfPBzh6iubxsGrfdnxB7zg8Ml4qTommgEf7xF51mnoOevDo6PjMjenEixlbTgAZ1/eFrwS
cKv/3i7WW+ePUbEJ1OeUVj/8E0n74/LX7K00lr2nYhzlMU0Y+setXtYq8fla9BFJFI/sbH2Vhy5O
DAqEuhd5dBbI7RIsjx7OtHQLfIW0n9mweRWcDj76KFgiiFZIyQuzJ/DPg534uf0FsF2VWwD9KsYO
ff7zp6n6pA61glPwDArueepvf0OOlFkNMFrTgVjM2q/e8cWMnUD3y5zuvjtnWqatzFzBhyACN1/r
q2tsWw+bcJGsCjoLTqwf8Rz8I/1hgBUiO/VAHiGxrOlIV7QFYKXtCxDuT+dDP26EJL1run89PcMq
IAWZZVf4g1k1Q1/ebCXER0iGjefNMrc7LaV8t4MQFdBrtX658fBqfDMLiy5RY4NuwJlOToHG/BaY
kKPQ/8k2OvbdIOyHNcwvwGtWMNASRjMc46X9OMTix2VA0FI6TgZH1pLSRGaFox+iAb/bsh4UiK1b
LP0Nb8dY1EbAF31/qQr3z3V+qOeXSh+zxHYgXWBjnZcTLoz0lS9ZFVe0uxWcgdnCn/rwaRHAKPLN
kqc8iOl6se61A5dx2WWwSysKlnGZEzwTF7xFRrNXUHK7ozSlpW2IcvykBMt0Pv946fjaQ61xE7OQ
2OZiIZvzsIaN8JCyCbVnFhcUs0j781Wp5qyIJHbCvuoT7xAkQQFsUGppwmXlDGmp8knowvtMAgE5
ZFYAnbQcwKC9/qKZai4+wQayeY1u7gSwWvoF1UZMhOfJbe+FYBUbvxYmMNtAxcI6xY9mEj33VjYT
dzG9Y3qnjjmTZmyS7kopKvUBsCLWadLIFioVdWqzrebDhyhp6fnwh6AV7gHyj3dZHQ8roNWBYo0L
5l6KcskOQmJ4wz6VCRc9kboNo5m7G+l/3O6uYZ0WpQhPHAyJ229RmsuHQXWGwOZxaRVwj3KuEtGK
NbzRe1H6LRqIV3q8o1gCEMNJ/Bhg+vv6ovDOiqId6vzPPs7jVyCH3YVxWOtwiF/egtK1LhY5Dc4o
4L3IsnzZWCeWGnzSQ7DbcLXhyUgtS4wwA6M0FI3uX1Zmo8LHpUG4KfX+4KUWqfPsKovBIaumya3D
gEpadNKRgHKUlzVxYKVvWr8A5RnuAHSXoWJSC0CJ+nWW/3VpL5k9zwV60GrvbXu+6/jtxpfUoyhP
8xXeQYLGDsvFPu6gt1blOfJB6wB7f4oSCJxgV+2wejKqM0d/6C1Ibzu0BLUqwGgVG+ZzccCVQKFC
KJI0bos5BSkMIz1yoOuL391ATf3Pl3KPCRvhsuGdmJhfBqAOLi78DhkgZcbi7Q3HfFoQp2KF6yBR
Jk6sPcCXDLWA98uYwU+jzrI0+mSdiLe+VXH1XbBix9/qzwXcjTvSLQH0bbjlFx31WttdWAD/tIUM
3Za7Q5mNVl6GMIQ6jsNw72gUq49RhObijzZj0+0j2qEOMfT6twS5tft+0yII7QiDLQ7mJZum5h42
7mA0+p0rqRfo8sDs+0ir0qD1mqtRtSD+SYqY2dEl21ukdNZ1sBdC0PRFAD7UzwY8kwqeh+/NeIIk
SmTdg9DF5C4FE64DrTawf+/lthwxdGKZhN5AK+R84ibKfzec52VGuWzDN89xb7pUbpG1dB4jrsn9
QIbftXMvL7vQIzZz1hoptTF+Hb1T1KErWDVtYXHXpARTKTosbIWLFuW2uoMNqgVPhJFDiLaMk6R1
CgAETfqx8SeMpYDTicNBMWa0jyRmxCFJnGRYqncUFDBPYcBZPw2DhTWK7dLdOdsIVwf19szGcPfZ
fz597AtxYeIthMg4iCKc8mHOcXlIE2ebM0QespIWQnMkxM5XG/S3+k8mwLC1/JAdxI6ycPKSRYmy
oYxTazrWm/973bWQXXc160phreznIhqwcoshsx1OZ7KnrwFo0NBLoCem0KnkNnXtYKZjGnEeFOYK
Vjub00qL/c9AL90hciyElpwxLg1pThgb/q05RCN8gAdW89/Xye1N+q3lsvamvKzcts7YsBzhHBR1
M5Vi95NsvaLuU2CHvliYxg0Mb95iAAyiG5ErGNt7nv6edI9q/N8WIDUVOiV/dQp9UPT2pPeoThdY
mpDJELkbVEiu4BewqeJoPFidmqJ4ectpgyr6pJVDHVz6tMT0WfnRS6tDmfl5h8vRfIfrICqLVz2F
mvCiVhZKchmi4k/c0DCiVj+tplpSZHtINYEElnt0l1A7mwso1ph4GtWA+T+/reouqKO1DizOrfIM
X67igzRXl3OFBoFzL5+FbVYinspEIN8DnKmyetklzZ0nEV3PZCxf7J7mhA+pQf6DrSzxIdccBYPS
aiNThezoVyGh5lD8l74Iqk3pY71rYDMOtaWSDfj1MsfVTtjByI6Slftg7eLppQU515h8xZEVBmoD
c0Yh7wQIkjJTWZhGuOU+qgRmCaKw0mQl98RVR8LG9ctonQUMrevIR//ONbLVAGB6hQsKq1uiLmnY
0ykc6/6e5ISgSPfuNsCwx3dMAFW3OvUnDMnVYHeudvFWCgNg/A/js4DXgRVwasE+Thk8Hzn3JFj5
zvs3vKMYCGXIunRntXYF0s3H6mPytVtn9aNCNRMWe5xyguRuKBvUX7cT9BvmUTpfpZFmE/DeIHFj
INIWSEqpoqJHW/y8lLyLjd9mvbPAr52vqbFkR7rzl2KKbG97559Es/sCUqGA9B00bzpPj+Fdtr1k
VaYRM6j9lDNQfIvhCO8JymXbPSKf/PLhnAZZhUxJuoQigjT1z4BGUbjlHEhDxNsGLDDWcRdBOUgi
UTs7T+sGAZUN+IjjjtGYxfEQHnbRNrPnBnG+mJMw1oYIxKOfeBsMbgIVh5dTH2aVMqxp/WESSFpL
FLp3CgrfgUp2IktuN8Y2tZsz/rXYeyEDUVcpfxCOWGOhs0krXnsGV7BNsrjUp4rkgOIxvIihLAQ2
gfMFtANt5FQ7wmwn374OwEJIsjISdjD+F008BGhXIZNX2Xvx7NoB38r92L7KyljUjhFgiuuptxZj
qZLCOqT0us3v5y/5YJiBgKhtMNotdOw3w9BYnD0pdsJOPEUsH09j5Rm9PrFclihPHt5tyXKtpxZA
cebVUndoY6uduOI4/VDcrNWCxiaRTPfoADVcuC46mnLhA1y3n5Rio0x7q6DGJs2t4ERdfg9IhwoO
r97JkDqn7y6W+AIMTvWGj3JYWQS5Mx7AC83KSCCLsbWC585Jp7/l0TqXRRqN06x3U0U89qZzVSpF
TR41cmo26ELc928RsYUHIFmZjnNkYbtuvC9UrTlhwbHR5eMlQHJrrKjXf4HSvh+CvP9heD6thbob
ret8oebcY7K5KTFeGuObTNszdtcAnJKq11C/PINM982ZzZ0Kg9Qzl0XgtuUx35U9gD6WVa+uNy/G
U42uCSyH/Lnm3fPnoU0mqFrItLs51gOv6MZHVSZZJTswFwONyIa7aiPpo4l89aexaKEJDVnGIsk+
F5eIELZ/nvN2hPPI/czLDbO9TlXqYpcD382GKIMsEtdMdRQZjQYjq3fHuM8nL3fnvjsg4TNmaYX7
a1cSkatxA6y9Sbn5xriJrip1MZC7w92iMiv7X0yyWwEzVR6PsISDBKSGuXQuasrCvMMyv1VGnhhI
ry3X+iz6ecWPptQ86RvMt9GO8PqF+i1gWDvkSxgcUAf5of+bKdHpmeruucWwQooczzH9eR+FenU3
9fLIJgS83p++X0x+bovXTyf1DHV9gFEaLTRS/2lF5gppbW0JD46sQ8cbUWL0kwL4w75IGDdS7sDM
pqsVSRWwocW4NPeK9pKpI2UWCi2jrvTNmGe6pErrMJ8+R3tOsuJ4zX5EycWfS/O66/mRx/wNO05O
IpbIAtDn6nZEO2spqIQx7UiU//K/xMguqvXeFXh8jDz7EiC2EFxZfzU9udH/0+HRiz3MRGuNsgUZ
qLxDgpONGVhQMhqdLYapMIfqNThT5Yz0MvQ1AwftGzlOsrjHV9j/a45tyit8t/vggb0ag+r1+24l
IlJjfX3WiOXCmFtKW3bFUo7ijv9Ts6cqzgqorleL36WkmYnOY9q3v0eeu9Y8PgCsrT5ouHoekecH
2YBq3ZCaMySyNwNh+mZ+SOA7Mf2MtB4W9+T4RiD9rthYN3QJt5II5H5nBJ0B3z1PT/aQIidf8f4X
lZvr1oQQdZpPKIV6W60JBtnPHkNTRvqh/36FHUPBlqfnIavO+Go5hkAqg/NuhS+MnTeN+eoSA9vf
IoFkh1IDbpuNrO7aGC7gBlfrqA309MifkVuLb4u6eCg+d/WflnMd3myLKkFmQogbNxmKHvxJ6Mow
g26RJQor018Jnu/fDEgNJs1dN3GET6Up57IsY+MwWUD6wFi7NiZ0iVIFxVlcNWXswv7/I6QL4Gh7
yO458zCmq4p0LM2ttRQCe+HUkhDrUzveYHd4fDx/VO3zJSVkvnOXWk8oPE5fLQjMPHOWUHYUYA7w
GSoE+qsSvdoCawB0ENyqn0I8Rjz0avu/sDUd40xTroPm39T6ouobXvgfCyxYN1H6+3TieIHe5vla
OZ2a2eF/IK6LAhi+Ml0+CMeT6j9NUKXYm3afDNULJ77kIvUvIoco4hDoura1c+PfjYhDWGaYzmPG
W7zT/wLb0ozkbodW/ZUhA8kJvk1iB0CJyqHJXOfe1rJC0vBVuBIpxjBfOCjplKqJ1lkxlB9/Jfsi
oLpGNyWNJRBSinJieVFAn5MeEhFgcbKjr+uQsL7TgjJJl+CtUtMXcBSuHxgpFTe+rX1xQXDc7/JY
ZBqIeOpvDpRZpDaro19ZXq6cSpWMsPQDaLZMJp/ulF2viWreYn1wpREY2qvsi/ina6K9J5In1IAK
f2NfGWb/jwLLzJq2c0PnF0uiykC2UkjKrihDl9liEtn6DL7qr1AuwZ9xOCaUlCcSOXecZy7FH4kc
Dx8Zv9Ij/+Cazqv3HTO/3lfZAhRcXixOnieo7Awj/jglCGgh+iKK7FEQZ4Myo7u7khdVpwtnnHoH
o75d3ApV66tarDym+edjnAEgINcQh67lLQszioc7hHKn/y30mjjVcEMTDGtOSW4IdNpbiwb3yqwA
1alAIAreY6Md+RIyMSBnS7HgTcd4rOoGuX71ZPhZck0i/m9BZ8gEl6r85xNjD0BVl8GTbtgZwzny
K64KUv5LTPue+eHQxWGcZzgWKpoFnkWNc1CD/B7QHLXOVIU3iWFD0n2vgwwgko0FMh2zDZ8Scy2N
+Sc/G0peD90rWAMGXzzdA8RuSQi85+wptThV0aSIqQdpRuSRggEmcyaHeDw0CbvecHQ1AterXAyI
DowiERBNWXPXaCh5ujR4Peo8PS7cWxhIYX281T9wp8p3LbFaXO6E9QmSVeyeK/+c1Yvwg9XWU2oI
xGrL+sgiW2NFBI+I5jHAiDveLk5oeG2s8PA6EBM0fCn5Ls2WDVVuXNfKsHjD0+tiflNNI4pn55gJ
/iEJvomuBHx2FyEnjSc8QoYVseHklS8V+/XRBtCW5qek1JQhQcNDv2joa5piKkes1egco8EephEW
UqKCNRe1ilLH9K5+PVXPSK1i5wvf5qeKD5C3jiiHgSWz7V6YFsmzhiZdDaD/1xdw9m3QDTsfgSYQ
ilVRf87YroVSK9sBmjkwCFGGi4FxlxIXCOUMe7ywy4TPvgpSmKERGlxTCNIrpzwnIGh589wYXfXG
oRbuN5zNwdE2tCPDK5xirpu+K6QFm0hUobzXPmBQuIFgiO+48LgoXVDKCsN8bvPB5+OIqxIiiD21
4ood7qWL7Jg0yTDCZ6g1dPTa9gGt2FF16o8YtOU3TJgCcOcyHOYod97uYpKkP48sH9sTFTmsjyn+
JUHlTjoRP+2P21hsfwElcbNCCjnWSNSIc17Y/tNMtqWPIzldwEK47D11AveWmPTWs+Ok6mWrYxaB
IjyawZaTOJPccKT7G8BpXExPbbWZAldV3ts0g2d4ya07HkTJ6tARS4fe2BQD5rTO+zx8tL18Z+Hi
H9xdtofttiut2WTYzwipdLz9PzTPLFzWjU55mYmgPGDrHQCdT4ql4A3HV398ftdgkfFdC95VEaRY
0qpSk/Gg7VfYLMADmP7LxX4jsjYzKaZo+nokYP4nW89l4trovicQf+M0gEFuOdbb0s9msd6ed9aO
mqeFp8/+/J1K9YSu/9M6/2kUrQZ5+1eYzXCfP+R2Xsp//xRyLBbJku4iAQHT5NpY0rce5gRcMKOT
REDt4AFKpwdV4KH44AU4w+oTca8UkEJdcFv7BmmD8Gx4dJ1/1DYzZ7mIw9LLS6ktdr8SHX6zwS1T
u6HduJ71LFoSeKui4fPczmrFKN9QRkjMNcCChzKIdb0hy3LZHWeMRSQf9A1/rEUjNMp1bt0xVoLW
2w2RuI9Xr5A4FRIr94oMamhyd2XF5JghwIKAQiBIHCvLgdgjTDxWykJCSvdt8Dr4D/1AdRDe4QKp
8+9CnBEBDVVOabVM0cyM4jXcH8DiEPfXR/Pcz3tYYLGE1CEKY9c4qY5mNkfHjjTglotGK2WNRnJo
HUID0YLHYtEIsWL8hOehLqsEYKRK3gVLpgwb7BfYPkVIjNncjB0SGTOJ/pxN7A6PRTOYg9ozwvm3
xhsc7H/Hbgz/NsS+ZjzDpFv/mb+offxzTzoxDjVfeDEnIaT3+nFBnvksA/pYX8I3BjBxmaocV+Xd
DWOde35cVH1nQ2UVtQkVuTwxZejhsdTodgE6IsHCiZE7MqJyFyRTxuK4n27bCy+K68nCb3BeLNAO
O4ZOd80XSsZiAWXD0gafmm4Zzx/sOgUOZ1R8+44YfU/mNW360Oc3CJp7EUjEQQua26h4grrbLaQn
7FNB9QpdNFMBVJBNn22Gvggwg+0OGiHXZ3pW5yBWE71oE5y4y8mHLzS/Uu0c6kp/kGxbLRRi3P79
Einjgxas0RxoC5QweRC9SBszLuT85Pq7ICPyUlam2gksRFl/+kyIGdAP56bgLkIp3sJEJulO8WgT
g6ll2uFjajmlaS4bGp2p8cowaQHEAtc/t/m33qThwgCs8cNZlmbY9mZcCkz57RwP8FWoaYQ0OwdT
uXxISn4L+ruQmb9BWsxIWqkPCON+ipCW8SMdUGHRosDTL1ndHjBdT4iwqO+KYYC8kXN3B1E9i+9T
j4gzrxkKOIBckJUHECPjWSu0r7evxWR94pEZtKdKiYXQzO9NwPmJy1i5HbXyOuB4VPGDkMHIOepR
t7D7th16/8o9E6tYk6bmekK5tepHCRMdnnG7zEf9TWvD6t3kB7G+lpwNtDFEdm0IK62eNXMy4vBI
6eNaJrP10VlUUSypmXdS5f/jY+jXraEAVQYF8uQT0E2je6/IINiN8+PsCEmexWX6amFgIpaLWYQr
lSQ0DcBcS2koqOtjRQWGviU014lOsGh3QoGlmtkAaMjuP1qJ/ckGwGoPIwSQG9eZmPe0KmdgWtt0
i6mYOP2Ik4aa+PCoPVrqEEVSuFJJtI5JfMzXHuXMjuV5go4tzawaNDSiZZQmi3kNPMvOiHqed2bK
ovD2mUgijnBHXRFVwCt3qcwCGlz7Eq2Pd7Uw6b7p6QOoXs8UGURmus/NMIbIQHXR7K9JzmOkI55b
IS18P1PCAtYTRLBVTBvdj1so6X+GtPVMjNZuC6M9E0Wdc+C8RZ8Wlsjoo+UTXMlh+Dk3ZFHI52Vp
TIh/dEBMpIrdD1vRM/8WASBBAbOfqxuOE9xv/SRKEIFi+x/kvvF3jfp4ss4ECeRXubw3ITnfi7bm
ZsiqlwTPhuElVrobsoxpP0JqI/ibfX9s0EQI5dbSQInKkOdzFhjPUctfQhEK7ltA59F8bSjysJjm
/C2GJShueyXep9XsNY5f8b+i3F4U16yKOhWlfgMtUoBOL5Yv3z53a6qbWuI1XVbzHmTlzIvqALer
hhHSVlp/6/9O2Hbv2tSLXc9YWqmY3rzsPjcaex3sqvFFhg0Zbg8dZFht969fZ7AZSAJgWhGUmoYA
KxLH7MEAs8kAqi1klHJLLXogGGZ9v+DSzRiuYlKb++KqYbe8ERrkYfE70i0NG7ZBcVRMmhi0kEnW
XgT1DnkO+FNV3YPtj3H/Q1/RWCIc3ZE4Kp/UWaHbYh/HY99aJNfiQ/Ia5WpCOpjok0KD4qXn0TP+
KYkq9+mbt5Sk1leBnPdDST2ebFUyDJEniwsD0ssH789r3DtlSjpFAESzNODiv0O0OO5aSfjb1ShP
NsNZ1hMTASqhMWa19edZl2/jE0ZW9UTUd9T1ZgAG434nZdbMfd6++rf/5W/SG4d218OT1XaZS+WM
elwHuxuCvHJpZDx47sKBjHCYibb6PImR6qsN0jGKw1ZxBNfez6NZydWHzFvPKU6P8Olho+Ht0oYy
x4WMxV02FOVoMA7TTkEDgvRBa5tKNibdJP9Le/i+qmNpoiQtKjM0ts9F1AFueQqTO1CllWR0DerI
NmnfeI0veDwZSJtXzKzYuKwXLYeOHDeHoevKm5EAfxNlCZhs5xwLaHT9u7mq02+k7uzIJ5JcdPaw
SZCkzXT5pLfWJg4bF3yu5+QLAaQ1beKxbYUWrwnk34jIcgH3AWslQOEf0WSkw6Kkv0M5d96SUk8R
mau6aaDjdzNYmlnmm6LiByS+ReMhJp5SyjFWxCOnBf93SUSOTFT5kOYVVnoFad1B2uIq/Hz/dgk+
emCItJPYsV04hpA2Nc0iF/7ODa7ZFmhpqFfK/4hG+1mGuzPuXSNA0Ll4RXPh0dMYPBkhUwFAXjL3
k4Y0OwJ63zWClXDSTBm2QyhTWawxLkR0LIwEd4TwS6xUwXrXZ2dh9nF2x386MGmQEZjhGiKyTGK8
5YhpZY/P5Br6Z7O5kY+K1by7/hPI6hU/jvzPkX9s806OKgljlve8lxVu5i/PtjRV1hiRvLIh0NPh
6HGE+dO/xv5OBFZHPOUTwN0LF8AU8+M+N33z19nHHbHbdMoHDe7cQs5f6BI4c1E8T6ZtNCaPfZQG
3IWBiotLi+65LN5WfXV5qoa0vxe6qYcgkGJLTf/Fenb0VCn6SM0kelKTYmGSe2NPV2G+UP7FTCdl
tTkdJpVFhYhkEICSX49lBHS/CxhFB7dsBM7NVBcI8XC8SeD0zE7OZbb4s+2bmD1zhqCgzONqIlwp
7K9uzhYWamI4J0YwDAxyLJ9Hcm9335kotsCjq4Xi8zcNKRgvXwWcevTv3r57zSo8anVNopVJ4f36
M/J5E9jpl5YTY/YG5hP2WOKEWns0UgisGlM1c+Ov/I8Cwt3gH7eArnjJi10ZqNrXNW72T8U9FraF
WD+cEhbX3Sz9mNQCUslP2YBrb3aBrQ3HWaYJ4WcIrArbB/oEzbnBRfpi59PHiXZRKzMZcAbnnNLA
GbwID5wBdWP6Wn2KgRs0oO/Bbl+d6SlKfhPCVPr/L7SZvAcq3Z6Flhaj3BNeQNQi4WQLvbxvBjWb
ph1bBLIOfC0idRyOoKch7/geiXjnPTau2AKRs3Nr8mtgMrr7+360UULjeNafO6ad2mL0OV176Kji
uYNyx2BPx3rC8rwgQ+gD92teDkgSO97/SqJBUsYVeONwwUwqLqk6jLeqE81FFCNFwOAYUtb8aZsY
zxPtx5yX06ZWAUIsi5LTcwG8DIluE0h6fwgWlsbI71L/lLqde1mTpArwA8GWglWvpI/Gnq5myjBG
NKcn8bgtlJgfT/v+qKLR55h8btZBuiayhPKyOu4ieo2RQCH1hdodr7E4wMC3tRx6nM9DQxj6nuEO
xe+6udG2Fmh0q1pjLA4hPanjw90POJLM+aGLf9oVDhV/rICeK4z8pW2UHbB7YapGP9mRvihGWZk/
rOJrk85NunGOggFHf6iOzG96qxFmGrdzdS67CW9Gcl9rRMjrHSwUxi0rJIHm6VYKtnwBu/Ljqs5e
4EmR9nXjVY8ESsgV7ODrWOBJKse5sgd+JScGni7VT8T02zz/DyjXs8M6Yc6txmUJVJdD9XH9zFU2
mkPDa31U/sImeAt54e7ir5e+2ttMD4TWqDtprE8xS5mslfL9KGHm7wdbzPdFbQBMA+vqBlGyuppr
JDLAfmOJltzMWIKt2F+O5z3eKs5mKDNB9sO35JQq1bxoocs3xEQIsMirg1WlzgFuFTe822OlMZ5M
jAJYsadCZ8Y2Il5Tgn8pFyKAFvEYZKP4KnHscKv23VWolQjql3W6KRrygZQoDTxpiyKsHbYkUkXw
Yja+qyqOIsll7L/o0O29YdTEmglluq5qpkTgrLlca3H96TnHVwyezBbzya02sxKlvQTX0Ww/cVsS
lbeZrdjl4r8M0vAoka4XMB2/xnzIzBUQFNCk0k4BW6RMvjsVPoSDOAoOTSU35l/Sc1+2L5nPjlVM
pe6jxL00ZF0Fmo4fH7AxLeJUuO7jMPtORRugplgABmYE91fioDrj1Py49nef0KHDPSgw7ftHWy7i
3up6TsUBXBMTim3oukJYwlIfTdiTRNaYPWTFyB5C6B6WhRA5JeFs5/olhBF7LazI1Xe4+MT6hF/Q
tyugIr+rhOV/djkjAuOO+1dBI8sHmNsERwCZEejijlUtRFhiNQ7QIQEq9rSoSxoP/5qDrukgEuOy
TNPOerGitI1WkxOF7M+sWMkvQg4TTwDo809EXI2xmHwsiRYpgYd8iUDVjy0wZUlZwMAXSmizyGw7
2n4cmU7vI66M4SK3BLh/M0gdSHMfr1lfaZUN4C9TM1DMe7fWTO77orLIZ10WUr2GPSoCfgr9o9Sx
jnpJaK9Of2godqb0fuYHRLvbP2/1kaD6G2fiZons/VujnGUMMWQ7LvAd8u5B+z2ijEsVOHQGzA/w
1zDtpGin10b1ILxERtMNiCUAYmM/n/lG7wHZz5Wy7rPDlzf9SkdzghPJVjSlJXExFa2TiLsJOx7y
EOtoeQnC5SuAr/tLEhHZwlsDGeidWdGkh+lQpd3soukPu+Jx5Q8c0Q+ttL4gLT6yRr5SPlJ9SbO7
VVt/x2BLz4a2Z0xeQZy0w1mm/0KYAT2sMaj0Xwc8ZZF1m3h8jeetRUTY5qGriMmixR4QOooEwdRv
+KmNZtrNSOls/WpQ2p4kNfijmAm51iEIHsgQ7pxV7vox9E5Lro3UeYMQrroVkJYBAxgIBK3YyKoH
0nBr2MaVq9nqLSFwOWtlm2F7qdJJVW2SYEOhxrbBy6XU4KnaCohq4Dz5PvhRhrIMzZHbfKNwMpB/
/uqUc22BxAqk+JQ3FaBzE9FJbdQo4qfMHQnXalRKPEw49mnIcJmWl100k4C8/jOr6EL8+LnDs0qp
DMcdu+50GNstuOLYx9SGptYkUuu/Lu4ir6EHFbSaI8UVONjaeFNkSkKKxi6zq4HQH8LIkJn3vXSb
KjDedKAmyw34/71EUdh3j6vASDqsUt3AHrN0QEh51WAHUCs5RtK78qXxG5KRBUP5nkdULNVtG+su
DljaYBmzAM33P5EhYOb3SRsslYpFLXyhJbN1brzZqXMnvR9lS9AwoYUO3yryIM59LuyTB5h4G5nX
VJezxzyhosNyZqhY51sC3OZ7TQb8x3k/CKUg0Jq2JoZwjHQXt+zQ8R2GM1V+lm+wypMWagLqi999
bhiYcXf2S5TMtwHu7QL915EJgMbYtfkqdXsNReJUtXO3vuYTmijIm8bmePGJ897H7wQ+iS4WLd6R
5HqfUN7lLW4b5eRId0IGbxd3vJo3iWoDlnQsmAouwhEFoQC1fucIpxCRypQn810/e0h97qBHsd4d
yE/ZB09aYFtOT7IW6PIkC8q3tgow03A/oKWbpXBA4X0KxR/ocfI3TFkS/MiijaoN7MmOBxIAKwdf
uJK/7t8KUKxk7Qnn+p8ePngAV8YxEWLz29pvksJEq6zqk5eFa7VAYx6u1JiKoXug+FtIZZNNvrjj
TBkVze4sRqnAkaA38GnTorIYRZSkgUJCgtECxmdYCcsP1XLydPZOgd2uuIYtZn3al1h8+FKB0EBG
7beBcl9YZCZrik7JkZE9SoVvacs9Yc5sortPqsC9PNoYsQChGHP/+xBkMeia+oTjvV7Z+3jf7+kN
zUqdtsZIflcbere1dUnDWr+2djXOhjNmMH3iUAAv7aRlOaFtc8g83zrRmOiHiOzFMDrgJw3aPgLh
ghF3DYavztwtjXG1wN1SOdB2JjZf7QZdPbROb72nt4gYvDGDHk95WBRE9cotrzIlp0iPfEN831eB
5+A20Y3XMSIE6ZV8oOAsAyzCWPpdBhW6F2wkuRYxIb+1QqwKcwnoXqDQ8p5VxrTCUe27rk+kMin9
LWl5PR0zyGTwfPW5z8T197OFTx6cAHneZZ+CWIKRL4MJ9wy5EDz4iF6cumU1Dd0pDQEf3Fb6JDf0
SsYCGBRVB8NZQQC3//oKFbpm0j65zEymdOTm/YyiCZ+/sgg8ObjATiHcckeH2jmMe/RE84bSbQyP
u+nbeWFf/K3p+6kj6DJ4z/iHEHo9BNB3i0PdsADEiH0UhxObG34ZGTtsZnIte7uOfrcyynp1YQNg
LWNaD8Vu8X5zMuNzBCLoOMWmVaivJhVR83almzqqaBqyvsb9IGjqoYMEeX3ZI6Z4jMJ5R4SPaDLa
soRv9RBDSsSG/kDC7cdl3lGxBBGHuulqpkCysYC5i+E4NULaSQUOkY0TEQBgCbs3l/OXIHOFabHr
e8+JCUbcE9+TxasWeEjHiC0kiAqZBIFuEGIVRycd+wE100xQrwQMXWi2qcwe40n/vG2m8hKC9cf+
wlQN/IL2PkyBSyEULJwa/iMFPdrSObyJsMd76UXizY9lnSFFdJqNFlj2IahEenxSxNuMRaznFPrS
skpvSeOKMhFT6GNd5kNQxsWPRKMohtPYm3bsVF3Rm+61lbZBl6GsSAtIfnQbNbUFFW4waDIV8RQe
t0/ARsqsVCBgH01kLc8nNR/zADKdgTuqt0p4rYkFoXdc67VQocakT5OKb+vVC/5Zw72hkiyNPZCJ
1uzlxGp3nB1iTu+cmwStt9IaSHn+0F9Jb9gKufUUr/u3lvLkrCAc2w/WlEg/M2yuInqh55YCY68p
PERfDHL6Lhh4ywFBknTxVH4spUj++rjfgUiRbtSFHGfGBOxMySFZawA1J4LKUpnmRpF+zS9pV4oh
2gs5VLyBDjSTcQzJoihgrM9+FN7nOieifT2uKzMG2yrhgtJokNVK3HKT5DwdHrdp8/Xj5pvTt/3E
7z40SToabq2ndKM5WVSnXwhr09Vv5dWyQ1VtAQrAGLOic8yjm/2DIrT7D3ijGhj0NgyuabAzoV7A
zmweClQ8xXRNus+VNN598V4O466TVGOcXKJeobF9Ad8/CSZuGdK34sBBWu9RLbjSNYxX9OkXMKeL
ohYZfMr/2PLXiaBcqVRxtpzEOw03U0U3YFOgYLdM4UQwSz5SEdzzFgtfiBD5rDDpTjE4OjlZlsU7
8PXh/tZL2D7DUk77/y3LurxVQdfLt/MrpoMJqsMsddAaDtNVd0p5MF52T6clCLNjZWbiQuOTI9O0
n2a5ELgRbdfTCQ0mlCD64XdrisfUcLE1tM3+3QK0dbolMqcszJH7ECNxsq2xDB+Pe5xDC8G2mO0L
4n4VZabDdqdD2cIbK0zqSsTAnKvBM9QKQcC5defKBIQD1fQqHvyZwDhaHlNSl3Y9SGXVal6X5Glf
hB+DnpVycwGKQVSQ4v2EVUBdls1pyWCe8l+WumVSI4qy5DUQvLkvclMENKnNuW+VYfyJRzwCCiE6
EPD2lkkTG4uiVWveXUDUxJduojr41KnJK3NEiktx3JqS9aztsl+zUAOn93ep9HyWcICp3youhO0k
zsWUMZHmzX/asw+O4eVSuUZm7iYAhruoDOP4vUGNUaOUHQdUZy20tTquJa0lHUhC42WaL5iFSP0h
r+Egq4hnc0qfGXvKRJTV4lCDoumKoqGdtT6M795TCqvwkyBsZR7mkTWmUgg7WcQSwwvaZGTufsyL
RJdBi0Rn4h10E86CMwc7K+LVX7GM9DoaTKURvhmRR2UhF8/JMMJVvA8Hc+RCZ1rXJi945AZcqwCo
j/Fc+seDGZ7qOxN1eRjOWAAsVh5aQwjED7JTotRWGdcGW/VX4ygI/g7hm3dRS/7f31bz8+lR6mG1
NG5v/M5kvkBrEhfCbaQYHW3pe4cpNcziA26627iKZnQIzpGbF8rxeCc1Z/RTkgHpmGVvAcrvYie5
U5PJgF7t9TDnbG6qAQv7hH4NISpHZ9rgIa7NzEbs1CCQOD55wtx/SEW/K6QUTD6nCilP4rSg7kpg
KhhLah3y3MpvgqgSITQ94vTC2+Ajt+ZSx78kokrllOE1uX5S8IrmeOO+yP7Ele92O+rO6gNJgNBp
ng0jBcadEhqI1tR+vnTxm7xZIb7qYrdVxzx+bhTlvrNo41rqiShSNldX9IHzmiNna3cKAYRA30m4
1X5hIisqRIPkQhURyC2gifdeuKuXgikHluARJMUaimypHyqg6c2i7BzhhezDnENAxL622Tlpz306
VhvHAIzuYIwQITL1PnSs6qQowtZGTTaUpb4P5Rd0jUMLdaeg1pvsOw3EJWnOdHHxLJA8tHpTeK3R
oRP/TBmXSN6eo4VnwlJyvxL1aK2dj+Yq+aDKRXMDIeuzk1WFDUhaUlaAUydACwQYt8c/rlqz84Nj
BT3zwo3jcCId7+QRJe6ugL+n4lSleKbBZ+WeRePpdiQl26Og0Nwx1xnNUUwZN8btF8m2FUWJflHg
HiquNQyTT3BfNKm6Iw0CYBDGmwJN4BHiqHVsuLkebo9TkHCN9ZEHPxHfylPS1VRG9L8q2hO22FsS
v47p7hHQkgMbf4XAqWL3Bl0LTEGjx5iKkEQzbUToLOBUnMc8VK2njTIaOmt3fqbOAcimP+8WE06B
vpRiANgnFmgdZXYG0b9G+rNcestTUrlB5NpXaaCy/bFj66omDo0G1G9tebflc2+XEm6YVC6bczbZ
cpw5RMicgL9ocU0h5ZgdFDDFbvQzQQHzS7R6krmGKqnt2iCtn/smyYOoywQu5mgTBI2GHsGQCj+A
wqkVTOog9x2U0OLHeB6KanEAw8OL90Yl7nC+HUTGL9Esng5IdWZlJ0ra/4XbCE/NHGKpMfZeWd8e
KCAjYmEo5SnkQ+nWKJ+sPueDDaxpbL4DRFYdFVWvlaEA9qcJfo9F2Scaw21hK4FAPQaJB/lirkl2
zHXq2CVVvA1oL25a9TVcO2rFRd/V9s/IuI8RNrpdgKu1Ou1zl5DC9u6ZVmA5I/HIr36uvEkMNAPD
voUCuDYVcF4xGqilGdlAAd3wunRgspCj912Y6qVpzaEFQxwhuBy/CKTR/J4Uij5+JtFaXwofvYjk
qD6rp3Di5HM9Ak700XStAaIokgQ5a5/rXyeLepF9SvQSodEeiPKggv0KQpV0ZrJVnQGaxfIzjh/O
cPjcBNTSzU4af+EcFoUEhyp1Rh8R4c16ETs3RpfzdAEXJbD1Hs1rQnDl0By+b9Yd4e85nKMzTcgy
FAP+Km3FDZp3KKE5rmzLvL73UOflW2+PpH6tWo0UO/Shg2Dwbu3/3oaLj3AKh4tc9RYXJ/eJUvuh
6EthqdxAgJmnm63ac/ivJuWsYatO8xrpdpaHLqHo+2fXZqVneu36xVo/xnGd2wWZq+xQ8wehcw9m
Pt0AVoLXKV/10Ei2SBM6CC8s7NMRtYEa8OhvFfhNv9ITScOZgTyg2kMTiQUKY3n7KCBDqA7ZyRCS
k5ctgxOqi241ML3XKRDbFVtN7YvjekBX15jmGAXHY3kj8zOBK8TF3Riap0w5XXnPuRm/QBxTvlkL
NvaCzTDqupIjnCadTAn97LsCw4IZC1RGlo2YJDyIMWXKvqTmiRfsxxq63g0RgoHYhiD8RR7NMoyK
X2Pe0SNhF9BnGrmAX2Wcv3N/e8iTSUCXdtziipJfH5/UhVr+I94zjTD5p7A/NBmmfvNGVIqAj3W9
9BVhuoM7WErEOH5XVKLdxRBnqFhB7cuJWVFP/IdZFffgbdLWMcRfRrD4ZQxAnMlSkYis2tGdSiwE
CxTe0QBkcWtVLB3LW/fdLYq5tyKA4DU+ylv5UmX2UMmMn4hvLaGRRWY8twLvPQ73tn0PyNQSkARg
hLY76cUEpRWoTlgZQxfUjjdYX/TJtq4/1uwan7wqTRw/0O3ZKsL6SgvJH3rcH0SIQbWTgK8K76T7
sDhLGDjmqn2bFLHHLGPrcHG/y6hFYhGVPTVXFf4BL4Q8Zz6ti5Dppvs+ulejMaCDAwTjTCOLmPtf
5US0/i5mzC5CkDBkaJFszV7EqL28u9Ni27J2AE2mubLYYHBt8L3csLnkFsWoriBGkDizJz1lFyZm
oh3Cp5H+qV6j+5d0nHN6kaaWnw9Rbii1aDEFBMutUGdK5+3ot6sGye/l968deF+CMMnLqlvh7WXr
oDutSbyI4ZXlvWLb5aCf8yXbdPtB+eTjBiNZKp62Ui6ZHscqt8pL3xJ13AtQ6zQCj3kpeixyNDaq
yhC4GNxuZtatdTPCK/eyyo/rwrO+gNgXYO33n7LiTYFZVw6qnxq0hK8OXPOPcVraYioCK1T8Dwvj
wrrYGJYyB7Ji8YHCf25qsb+E7H+Rjy3phfopICvxAxkMkvtlBVcne6EFmkpcbkvCY1Bh6MsVvak8
YhfvUDk2V6r+AgJTlVxO1dHLB2x613q8Q8GOLk0tCvSmpqN4jdiY6lzdQW8CqeWumg4DE6+A2Prk
MZBgq9qIKt1RDJaWMSGBmFKUV+nGoknHoroRxHc5gLPtZE9eh4GffihnOjueYnEtHl/hun2o61zp
LoJ0msJxdDM9vJR3Mm6v+wuOVakPWPL9KJVZj3WSbk4gBLPUbl5FUcpJbEy57tN5AkoEO56r2Nrv
EItC2sQYGX+zH3HNVdRaH+HUX1REO/BHp10aVYVjwpb/QoNCz9fdlJT0+jyxQn+AurN5oe/hZZz1
tIHVsO9xhx63KOZ3Hz7tv3sBsSlWy+ZmSPE0MLiQyTmFt/kGB+S+f1G2FOeBkQ3tfarpBG0+Ngjm
YLmpFmbJV2BqtxMeHCmd5ehenXIgq8pFAaltHSsiM+TDNfjuWxZF5qY/K57H5XyB5ZX0wOH4FtUO
+OAl+FNBdmdCV/bEmI9T+I1ufU3/zBU5ATdz5V3rM/dIyvcHzTL1W/UFoPNZ5VTGDPRIEBKjJh+A
T/q41Pv60lCDiG688lFeTNJMVTXfbdtNu4V7D3wICruJAKSJuIExMougBkYpQw/Hsby029ObSjBG
3tilvyzsB8Fyx7GsA2BaOqHrBolR/iRffS6m9QshfMy19XsqgxSmumXW0+AcxqO+ZowT3EavuM3v
GoxF2w9d/Qigfwt55iQnCGzTQj2utkfimGKUZO6K8sgaKQmnGHMyL+LMxOVcAXSHXdKookQvL4oM
CDOoYgiSMfmKh5zr11ROx2H69n3FIO5XklaeKM7TQfBPakPVq9zXp3pwNcHGtxUQ+hwiGxlEG5yv
S6V8+SMhYFfebYaTUBa0jEUz27bkFroqr5utZqdl/7VC21vt6M1lIH2hWeRkVuCEeW9zDHd4NruR
vcyziJFOBcebm01/DGg0OtmLhV2AvI2l75DgtGJnqL9r1s+ZpCLJxhoUEApQfI6xxpmxlTZSbtPi
VZroGGz3Snym/yKIBVayN3OW/gJuXa34zR3I2BcAANqiEATT28ZkcRYxJe2T2rm9emDaztSp/c9C
7FHuBjoltTou/54ReuIuPSn8GR7WLnJJoHbxwhoSfOd+rKbzhfrq4Mf2L13hIoLYAeotPo8tZB5x
7ttSchLOWmviHQYIme9kiBAbvtogosvKbjVPJXTzxLS50bZ02NKEceGFPUGKe25sUZDxIkGY5f8Y
oDxLbuNlDbz2Y/ofdUsC3k4Z3aBdq+ooHMSzw2ATbBBq7MC9YfIXWFddaLZnUMqlZUgc/3U8VU8o
vlcLsfKmesDo+Z2K5STYA3IIN0HJEZvngVR6NBATs1txNJ420XTg124tGvur76Rs4nfUGrra2B28
r9vNDXClPwrwkarJbYNdc7QzDsB+lNdMfq2X8reQCUkvfJ6o18yQigGop3vt3U3Rfyv2X1QwJBl3
DduB7BIpNP7p0xXJdvKdjKaEqq6T4SGFfE3JRJTJtDpZBdT3Po+V1irOzq2HeTkcCicii3/B4tDV
S2j7PDYLrq9cjSdR9nxfNQYmFmfyzYy1BfDherihKzOvtt3KTNLLykMBnsZLBYW239+fzxICbSYr
W29yLD3WKyZi32Ka+coVk2l5aINYFpn+N5JvypZjNfQiAVwsEszn2Rsbpfb1u3BRhBfitFLDVqA3
IBhKoSTKU7Mh+xLmRmnROEhuNWazA4ui2B7s6yZm94Ps8JJf25DDeICa6kEurK5Qz/eQcqULcoH/
MlxA0237QSDuTsSrfXMeNoTlr1e7OhjwOTu2D+dVerHJ8+Y4Kc2AHhdURir79b2/gN3nNbAZZfVY
rYwVbrGIGTljbC9ojxNeCorOUw4bpjBoDpWGCCdD5PNc/+chqZidnuDrl+OKCvoxL5i89m0b6AwK
S9TyHR//wT9rwOky8e+DaktugAf5cYZZMY8+iwft9WluWbuilPrSJbgIK6CrC35X0XjMhAJSKIJQ
IodlY+D4PNF8doZcgvt/STEVllj7j3Nzrio/fGUtiXRXaIhLSkr4ePgrekLqSgzZVVCc80Dg+wcm
cvAw+XsBuF8b9LUHGUZmHQMdQryAPNokf9Wejy5Q2IzCtPIHqbsauIp154RYu4duHytAzm4TEdMo
ox4dFAy3L1ftUM98Bm3CmIxwVjAL/DQeH73uYRjwyjbi5He6nIkAbaJa3GaN2anV7t86BC3WuyUX
O1gnrvnd5js6MX9QV+nd4DDNXUTbZlrDoowDZBaf5J5EQkLgzLtwRu2+0+vHCNOYUhwhoVZ4jpU7
dBP8+/oxQiqGEovlduyQjdK+Mvo85qopFdPfhyKlxm3X8F0NFl0wZGCngARooqSwyKLOGC15VC8c
CbzwHggnhLyjV43O+pK7peQUmjYD2F3S99G84vikKNX8H+Z31j2mNpB6S6TyDJIESTH48laTQ9P1
eNdzzy1BHnJzoMzLpDS0BNzs7PKKHbHXwdXifS6xJ38/6HqAiiVNQiuvX7FgISjPLWEJa/41HjXL
olpBuvb4hze2HX2rusVaMyJeSdIOvbo7gAYomcxNSS7Qhi3DbX1QQcde7WmCt4as/gTrajPUJQ+u
KZXFY142LSLaMuEBhpluy15mQp8snjpLR06SOwJMIMjxfMi/jIQzTtsZkEYsnTSTKy8cy6JyW41U
U/F75otjb708Q7yJdYny9GExAXwpdea/H7/AKgXlhAMxycmzQW5kzYmO8erPOgr7MO+Io0xyRDHs
GqdoW50tDxa2Kyc3EMZo+NqQ9/ky4Nh4x9PquTjXQ1cNDOb+XV6GBnOuJ4cuusw/6tsn9DsQSpr/
d7QonzaJ2pv4rUwc1W2jbZrJjgltjvMt+M/oZSciE4ZXuw3cjioOrN56z92Xpf2glWqfihOzjLmG
JHcW7Pe6pQ2Is3eEeqw54OusRYIRxEfLaXT4fu8RiP+PSSOlKQ0CNB+UQq0adZWeV+pLA+1cvUZP
qsgWR0dSAfsWxlPtZEAO5tb7ItkC1Z1nl3CcU1OoL4pImcXFdSzr9pWO7uyjlURZxaVlQr1zenJX
Qz1YDCV2DDM781f00lvJx0RCacZPIk2eq0bkneVxsIWulSz8bSl7hNKJgQu416OJ171+X/XunW1l
bgfiNhtodM8B1fymRidu+PAD6wOEYBbCLdUzc3zYqeaw4/kvnH55pqGaGICiM1PObwYPWA4ORBiu
1Ji7t9VvmX+Y9bi4D6VGd3rQSb61QXuRLCNR3+FcuC/LdAUV7QIzbAMGWHDGmeQZdTwz4c4fjEdP
/8Wv8RiVn0UxvlsTJxOjHl+NBvU0QAm02uM0zmGTO+1tk/dXUNZ0uaWcjhTxpIo8V1pYf4MZ7mrB
YzZkZul04XT4VZVg5XOHKqKh9XT7+4CR4oXuIjQt7/6CTQ1ClWGTJD/pepibzMINLB5EvPbULvH8
7368I9bEzYr/APZr1A/w59kL8FRnXB1O3aHcaMf/3hiZc6Jke1fEbqhI6iFJgEsw3Vx08kiobQcW
Ke0Ry+VO0/WggpU73ovgFjvZHYfyO9qR84NJWrO+7X2E93W/dytGFlSt/4IHMFC85z9vB+fMElhu
1evptuaq9vUdUsAOIvvDP0CLFQ8n4n1EdmuXZuUxonqUjIJ738EixgiL7eqkuZ0UjZBAPYOy05no
BmzmB/7aT8VzmBbyvkGYfte37+OGLfDXNVp7vnxiuPaLwInljenIR1WXD4FkbuuSjbYS41WiFWn9
t3wB7kXTvpE9UwShNw6oi9EBWSlni/xd+w6Wy3lFyhrw8bQQMvEGnCos89DvRoLDepgKvcuavaL6
bk1fV4vJVrLLGzYb0GlavVsY3hEnQSWxEPxdURjEFEoOuhw5v0pOE9d/Vrqgz/j9W7Lsdp/MSn3p
mc/s5bbv9GTv3/h2naleKwQV5AVabU6hUDA0PTXf+M6Kbj9bPRxcPGg7AhobAYczksR4pTNZkNGO
1gdloYxxbWerK4hg13hzO79A1/6ctNExM8M5WIN751AXoSAoVdkJrSCnyC8EF3+kMLkirdgpXEWS
FZQFVEKkq++kNg60tYJT0csmXDQOkkfpmA0oM5m3I3OGvclu8htOwL+gXlO6XZpdHpsimvdpnU3I
WRH0FFLivN1TtA7dLSBNZW1uwLVfxoerScpRh14DLlCo2vEelejJKNNd+FWDxajFAi3XvYC3xkFN
LS9zAh5R6Fx+GrdT/a16nSACgddf517yR3Tjk8zM7xoJzT7LsmDWAhcCPFp5jHOHdSdhHKwAYt/Z
Yu50p/N4qDGyC9OhXpqe4NRCVD52ETHFl0fHSxQv0aXS4/hoeWy99NVXkCLzNQxTFZ7jwiEvm4Aj
3UMAncGqRK+Uqpv9wQqWkq0TrWNKkZ2iXmDwI8rUD/lG4a8+o9YL0WrdhvA2PKCh0M87HPxZ5qE+
YbBS6p5MI2w0QqeKlvunNQqBWiao0T6kg6FBnNfhSh2kLMSAUI+JZq7NTQMRY+x4+vF1Qo8aQkRq
JAdCRXilerS+rNAMdO95gdmTLsa+CB4+oMDojAZOZggqYsG4sCHEGfHVabPE7s6p4ZVVZZZqI6yL
fyHpVTEX1MDgVzsJ435Y1dcDt230tRgQzNfVvPu0pfvRHFRJIQnxNQzR45wBTBSzwS2x3qzXy/Fi
mvmLJqOC9hsQtXO3cn2jNDdNKZHR6/lWCadWyou9C0SbEk9cYJO30vOzZusaHOZB8xk/RXe3zPTE
a6z8jUz4lLRFu0Nv4VqCOR6ST2bKIl6T933kLFaWWgrwZzXaeoIB50pRgjMYYpnlm42d4+k6igH4
fxJco4k/EpOHyAZmI8qoqkve36Noi1fRdf5W59n/VAs/TDhQsPzGEaQezdA64ul7HdLQiNndDyTo
5Ag+1K3Hq2UlGGQi2v6yAiu6zKZnluwl+vt8wHbg/RYuQIb6nJfA08fz8Gp/7zZsrbw6obkf2+cM
ONqNMFDdfuEKOjmZl3ec5rfZ+lOTXLbRzHSFw+Knh6Igh/h2gH0fD6B25wTE24B8J41Bhsk+W1ef
NOazdPQf5rRK6MLra9LguCRdlG+VUn11wSYd093m8OPBCn+P6x27/mN1mBv/PoigDyNqIal53VKF
wkmEFf5wChGSIWvD6R0THJ3G2+eSSwfEduS65MLOAH6x1V5d45Wcsbn/qUE8jz+gyM5FqZbo4eFq
jOZxt/QUC7s8FkkCHD4Xhqp7U6kwxIAWFfzMbbzIa/UAzhXkEpSDCxPlVUUVinB/754OnI0tIKnT
K9m5ZlgMrnbYHxuzdsxcFdOYletawpb2tG8FIAvxbWGMZZr+22UAhwZqLx8RAB4wFGcYG0GCSt/L
F9gei91Gwt5YaABL8swHiItK+ke4A3LChEtEN3nhbuBHXxjdVPFzbje3vW/nfCjaYVWgiZ0LQH9Z
oAROO55I/x7p1hJkezYCeiHJLqsROMCuRy1R0iv25Rj+NnEdW7k+6i5//Gayo+6KdjX0+/O8mIPV
z8T7yFrfAFAvo24+hDVUfuTmvQsI+v2jD3HGiYr6eR7eiYDjijYcZRuogDcujNpLFE1H9R7Qym5Q
V60TpH16jTx38+i7AVpXaY1nrijmlrbug7mQQfZAYMUA6czIVTko0VXZHJ9wTi9SwMzKbwMVsDhO
DJfR5o5Sta2cX9TStqffPq17+MU5VWz49uf03cSSgUUYdOWRjOxb2BvsrsmQHisfilESp3Ece4Ka
n0rb4xXLmT0PAOS5aP6nDJQcaM6RUSfSkdkeYeXMpvQqc9h6R32/lmeEYrXo/kt5zjemyzSypzw8
fR5GzpIvBGErNDl1D+T+fkpTfWyldHaQrBBhhGRMDMt3V5Znl5hcvNEkyJ9F6qLiI/wXiGiGrSoI
ipVufXZqmFnNdZ05nsjTQGNce/Zb8ta81U3nDf57vbzeEsh2ZvjNkjALr8loEItuh9AckPHdDr7P
95UWYLuSKPk+FIUWxsSIw3Rzbwr7uSOstdBxc5MfUr1R8gYTRuZoEsLd6Qe/KQJmgq2i5xzaYOPQ
RWohrdAH3J+meKX8wLNJenI3jwR/XkNK2esr1svOIBPZ/G80XlhvqyAmS3zKlaIHG5UIq9+f4oA7
F2kVjqeDcON29XAzO7yMJoYHPO1knU5igJByoJ3t5D0MExIOGjHZkVoNKQRaTKjzBRWY4Sp2jsOo
XG0/EMCt0UudLzEdOpXKVAmxBJ575OoZizYvhrq5QnPZ5XGKgyy7q4PpBq+HrEjW4jJLYwhqdDtO
BUmGiDRdB7OW6MU5RZJtB2yauqWDs+cEaQTRyyOBIuiKuUFX2+N6+JFKPlV6+hvqamhsSRNJxtue
smG05eb67tezwkRlsYJd7TLDMTUKJsfcOZGUQ5+9rOUpg8Jd33jrYBDiELUtnNk0l1Lf0AnPQ+mr
6N28s9JXeN/o6dtyuvvOVGPG8pHeAlryxcHPXsEtAsN6A3mLlrOh7+fePIhjuB8goxZrY3/95dTm
PggyN2WcTSVkc7siH2f9cI9OqH+BchXHQSbosv5k+G44Gdah84QECIeWtGbeZSVAU/ao2DoActW9
snLMsQX0SvURJwAOFck3MmfUVI0efnS9Dh3DyWFjUd5hofKW9Yz5TTy//+TmcVyfoj81Pigq+/cM
3gOjrq2NN6okIhQF7VunM7OiWsiOdYG0ffFn/tRt6W34bjiTCo4UwOCKnLuAq0BahiDRtKq/ILUy
9t46BEfai0aGMk2gJCcXLqEdgW33y/Ep3KVzvDoLL9A1VTdyPfDkkmwvKBuLnpK9TQWUV9b5J0qN
dwBD2goZ/hr7pnv9VSog1ypC5uo2XZD5uHdHtrjklQ6wGcVVXozMtt0leenNQSHD8yiXnzhfLD5R
pRmsZbEfBLNsnldWrFDpiL2tqHbQTKKLEX5O5c6LkE0FVQZ77wqNKDaj2MjHFWN4hWLPjT5t6Kpr
m4WAfRrOEIDwKqnAj4sKnioiKuY8mGiY84nYYv24UqdBA/l0ICWhOoA+z3er6y+Hp7ANVe3PGXGG
OcdVJZBUgqFGDbmgCDp0+98BbtCwJx2qCC2F8coBM7yB2hbSNXuV+8L8vyWgG4ez3F/tckspcIoy
H+02XKLRekggga0sMaeNyyTsPenxRUIxoz0jH9eH0sWUEl/HpWN1Im2Uo3r+RS4cJSca4KPkMqt+
uwdC/09PZ04z59PZwt2SVsnNlQe3Hwlj5i/lMr/LsSA0xmfF3krnvCjRTs//P64Zeg86Crc95BM0
JpGs//kQkbAaWf0YtKlZ7sMw3p9CM3wqS0N4fdj4vjWuLllz5clYnDHtb84rZLd3j647iYdv9Tzh
1AJXwgla0FwpJef9V0wIPhuCzMU2BopSy5oMX5TpI2Poo8NqDNV9i7yrC/EEjrP0XIJ6yuk/vLEf
aXGiYm9azbn9mNV1LlJP8qUr/QYw4s8I7lut3HwBMUfKR9zI+DW4naM5OGJhllbbTro2WAobsm1P
RgKa3er/d33Fw8IL9Zl7y0Euzf4FNVE2y1p2a0nx+TqTnjx+898TfYQW2NabkHfNIoth6YjQxvgU
s3HXwKzp4Ml9uOlkQLYGt4wP9u1xs0Af4JUBQgUuS7mkZnBr3Lf9rm4QfCRZ7UmbICV421mBnx+m
fmubNELFeUQdbmnc0hmtOSl9nsSt7u3+uxfyKgJsl7ZDAIL3eEz0IWG2mwzBqeVJeN/9dDxzjjIm
0tHcwHiGGQe9hpJRaLJfewEDZfH00o2NkNNyIdGq+U9bSiDT23dr7b1XKGsTyc9jkEN4m/uUVg9k
f3mYQyE9kVEux4defjsDF/1nW+5nuKgcZXSRZ2EW74cgdM5FqdroSPhflDnasfsI5Kln6y6q6xb/
lU1IYSnzpibxiRm3hwmhy7B1GouvaGdykAq7uLQIM2OAK7GnJtxe+bkLLuoA3APLJFSYK/OOQ1kN
vpWrfAOXbDXxfsxUgt+fLpuyZBVDjjEt9CbOf1JOZqfiPM5i+FOLfA2sA0fvPwY3StBfYGM0OMoL
F1UbHsIiJUM7qpvjVWONpOYizyCOSuw1RaHl5s240G3t3MQoRVT2qapkyNVBcRqaBQ2FKCX1xmM6
R8PTG+nYAn0O6OrpISJDp1+MVu5Mp1VsvF/njqFPJNPnKpX2OExLH+Pihnp6jv3zFSMGXMVKShV6
yt8DYgKj1k4FW/diUbZWHYgOvAhbp1NYS4uZN8djP2WQeMw4aKdME/g2Q7jAA6dTOfeDbKROMOCd
ovqR4gFlwEqh4i4WJJEEu1JZGx5oDpzGBaEE6QxwIhgSgx2TojNc7lEki07g0nQlO55OY1CuxYap
KbzxxEEoxpKUuihTXqNCHwHmfXNYO66yiPcenA8CuGQjgGtM2tL80MSzNsszTtbCgZVPGkofy6/S
g/CZiHsIKGYiNnEw8cyzKzHk5dbAeB87XDpwW9QzXKOTAXLxMuyZhlVnKcerWSrYF3YVDNVoMlb8
wkJhAtrb/Y0IfpiccYkF9fXrzq2UdK4Y9qDTm7TTN+pYf7up/N/mDCK4lP7am64ePPSj0K8kkowt
XwY0ZltNopXh5sSONoKo22ao+DK0ushFiC6jI5BHZzQO2capa6BqCm9rbK75k/xUklc+A7un69Nb
vJzS0l+7q5EHnGLvBb/BeIL/OnHp0ioQRHjVhJW5DCmEHKvr2xsjY5CtZrHcdUkN0IQ1QbLFTVNc
DveOkVEIGGUYczDFrEFTPbmtLfefClE11v+WLEjmHVWOwxQUif3nEpbKw3bAxcqo2m7qrd7YEF+I
cYL1SYsUJzkQsrI7bXKZHsspjft1S67+9sp4+mKJvxoebmv3aCKDvTIKwiLVuzsVDeU2PU9DAAj7
iAvFjs9H6oEECyX3iCi7rTLISovbJJ1RDH8bfPJPj+WKO7dzeq7HoDLmk/MvOGE8VbaoPiAY6Iu8
puP/rxZZf3CYBJZ/Trft5Db8C8Tp+dE24172r86ojSixpcR2PgZt8X817535h66Mc0ZxAtqacKZs
a7E1Og9aMOe/QK+kj3hJHWlOxzfFku25p1BW5l8IFxXDYY2J7Usp2TaMl5BAjqZzuCpkl85JbQ8L
4yOP57JOYRaGmYg3Op3xKhipJCEZCJfJ2dxgyi6rev/oSkaQS+E2USP8uZB7U79VDRxHEiUnrywr
femmRDoD/AVJ9GjaT95WiwkS0y5w982meW1INYH7XCt1OtK3aoOD1girSwIbYploFTz2G/v2DJQO
FVBZ78daTsYsWB+anbjn7pYs2b7jYaKCswWjCffdmxDRyXeCVUifmQA7AEx8m8tfWxP3KP9oRGUC
I+Lny5YzFW6qlt0Sl5t7FkFa8VkYRYPUGcksqSxIv7WvrvAQNZ9crhp/MzK6066+n3VqzMDvBb7S
QY6vht4dnVf+wkPdfvvuPaV4/V83vGTLLhnawrh5SuxIzDRhIwTP/sS0m1sNemDkqFVh9T15ogF8
jfEJydVO03onlcPYKlt0/ZGtF3Ons8NWdjev2pUb3fW24t+xHgmLLTge9m0sLSYe1Z2cqiu9Ft/f
di7egcsId7ZWinmxMM27pvpmenTrv5fkOGnrzXp0o5c7j0txiySPF3Df0WtpWv8J1LTuTBKZ7XTb
FUEHoblp8Ua2XRxcxesFHW3ujDbDHvy6C50ZccU6Xuzoput4IZ+7zhnjahAHiOuEknriwvMBIBgd
b1Yx9+dH8G1sFLlw992X12WokUPcZ1LoHur0I193/DqouBplZE4TP9PwJoS3lpdVRbm/oyzIQpcN
8lKaTvS5WQDhG3+fgO4jWDCsCjiuXPW47KGJFCF6iWpBeUcZJxbN3fNxjAp69W8YdwwBEq6Etr/A
lFomdRK1E05JPQXhdnA1bfit/AElnQWG6ISr8SbxS5IsrSr8Z/daazzwVzS7npuFqaPvmMuB81x8
X2LQbSSnUzCZDx8ViTJCoVJWuZFQc65UPxo9Rmfa6l7043v7KAXCSwBZWUSKYIQVz7TUyaFae+Lz
6SKSuEET7YRzJHrMnfFgXWvvptY+NHzgZcJWfXQLg3vAdQE2KcEHJ+za0YdLKX/BJ6sXb7q2K7Pl
SFEC61/DQd9wA045M4OgtyttDn1W64tGBKY68SDJ8/yjUoJ+9DwfvW8bXhoXKwJdlBTQpNenzWPt
ftLp3d+mwkVqhaaLE9bp8sUG0gRGYzKyoajEX7r4mkw5kQb5xHlXnbQfbSlAWruxp0HS6QtV9rYb
7I85cjU4h6WV5ZP2dzaPER+D74v3VJBSrkQLdamFhdMzwrHe/1Ste2MdzKnLV5maFS9ncQtaMLSG
BwMjxWImm/pzC7iFCsvTSKoulUYS4bOI8gEAkOAe/2GVc95/PoSgONJCWbZIsd8qpWteePHgr2+Y
Dn/9KaI3ToWQRChGn2HfnOQcHKFPSIRUm3Z55YmUAXyAWwzpll6YAA5C/GkOGtalVXJA+kUZE632
UoC+jhCSZH9A/fjsYNVGD+jEoSWKt9L+Nt4fomaPkasEVm06RP6T4i6+ceHS5sm1J+R/2lZhJ3Eu
gSRkMqxz+kiRz8So770ZlIE0WUPw6+zvrFYFJkPtOuz84SHlUcYXCypF8dZiN4EMi9davZREL2BW
FgAVUBfPR5WyTk9/qm73Ed0jBAlkZwgJhnc+MtA9PE91XLQgmyrKVO3SbyONCnzhsohns0jqRFa3
qeSuhukL2bObXS2+RWjDXF2Ym569W4L+jMmfukIFTKmrjjPaEzxNzub8viJk3DCsDo2O6tf+3nT0
1pPu6i6klRDGLnXklBmaB2i1e07oBopHpb8PpPUeUtuPPXyV4R4qpYLeICol/NqUJgUqdLVTIi0F
m7isXMzZWkOvD3QrzRxh3OjrWshBECS6krHFq5y+1o34gL1hTIsxYgoK73dpeLYb5qsyxvaNF4gu
/hy99teTTAGyKg8sE6WzaSZY7qQ6cB7UwAKq7G4mT0CpKHuhEykQ5cVm5X/Q1Gwxx+HShieRGXC0
Zpvi0OHu1uY4SYpgYarZpQbiccRgbFgETKRtDlns0VmuvhRWE9kiNl3OdttsK0gtJpyFUYylZQav
vfVM6W9T+CcmYS225H7ILCvJgr/rvtcVbcNBjXEtHLft+MKs1CNeZSsS5rQTmVlDJ/cO+tnJ4wz7
Lbh/4ZcJkKrXMTdqV8mKh0nkkYnxwd1hvO7NkKjKXBsqUPmokpRNZiRMALdHg6b5PGaIS/EB3XTW
6m85A8WAcFZM+XoVlRC4G+zY74hXKtgL0TAXX8rOWmylC8Yz9/2PMPkC7ttIqAwp8fga64lKvhuL
AxurU3lMlYFOttUXZBRepdNP7zmU9VGYxkKrfMUwhVaAYFjdqC+5stPiD/lMEGY41SnFnbP5Y3Bx
TNOKi64ZWSbTi1LyhvmAe8LTHyqYBkiUUagV1mQtlwpsKcVSEav8zuxR4qp8mFWVy47ihq4nfq9g
YEb1wN/tQSp+v9MsTTUxwNT+qJx4SaK34PUt1xP3ZqyvVOSCdO4nmPrjlL/K29Vv/A5G30eG4FtE
wiWRSx0/nv/kB8sOpUOsjsIswWA841E3fNnOlEOuryFxveNgSJL5RHRlSt0X/TXY7EDKGsWIWffB
zhYnC3hOzbI5plzbSKQpAaPMaGIqikUXzXQoQcv1RW6TFnfnhv3EVkR6vA6JVdxd9HNUjN7oNGjD
F+d1O2M3+yVewf3aDmo1Vu/Wli2x75jug0ptB7876I1WjC50u71YaDJH1CWWegGGaEhjeujKv48X
EFu4NK53VNc9DOW8Fu08ohMb40cNF9YiVnMcWVuowOh80qfqrYzryzA9ryVjpcki/a6h4YFAa4Nz
ZGTXvlARNkuXV3H3bigpyBRUWI0FgTtHcWVbXyeZc3CnOuR9fKY9YREhorNyuyN3rjker6r9lnL1
th+suQYzwJP77FO1VSS9suFqktbjOlRtKqSob40v/Z2Ns8Iy+ocsMN68AhLxQY7urAFG2KDWUQ+x
j+2R2R7z+65OT5s6MdRUbhTXbJcL8grssa+IZ+tZ76+Lrlg/YU1HqZtnSRpsUztLwKjKKFMtr0d5
pPcIpW4wGxE6qUhJu1KwoWEgHNgwAoZc4LlQ5xnGCkSbbQDqegVBZ6gwNP7b325E5oUVMm6Bq/M6
3NvwCK179xICOuxN+6+jmhqRIxxAe25IO1crAXo9UYBUccsheB1cIEuiBz9r5jM9hNBIX4y/5qPr
VjFmi/QbHvrPO24H0V0RLILQRXuvJU/4RUBPWimChnoa2OvxzyD9gxWoMeBzLi4DMZWSqORJ/xYo
B5bEYOFA2QqKMkBkZiUE9Kko5eztChmnUE1zL8eJkN+NfOBeOQOCD9gKnk3CSPWn76MlEH2xKJ6F
y/RVi7YFv58ht5eftktG+HW22qqSQL4Fa3psDvW/NioGktyvZhh6OTyiioD8VBcuD/4HDbclDNgr
zCv8VzlWM/UZDBo6scqCMe5lKx0/2G7smVtIdLbroWxuW3bnYSLtYYfC9QdNIXGY6sKjABQp28Rp
iyKSN2e8jR2oPvQysuDnNooyMibZ8Me47VrYkvFV2YGl2dKGJ50C5o1IG1aeOAr4PFddwJ2lCYgv
hp3tGUu5bMspekUOoU2map+kTo1A7wCUR2sVJHzwFI8LVrnyY7CCeSR36vGZHp1BjjcdyK0htxKf
+wSpL3rHLa4p/rf8nW2vmzM9kEjvJig6MYsXW1/+avAM6Xm2PCB5kg51C8wOBKzDvSztsQtjTIBb
PGscyGJ6SsUsh3HB2HEap+WrmPfKcdKKDrkPqv7tOEX/EMye3bMQv05nJ9DIi1ytBWo4vc4u31Z/
5XWl2OIRx8jIXS/O2JX63tWonqyGHfTwodADgopwNlTDpzqmK+wVEgK9db5rlTN0Au21OctVZ1FV
dcGYEOanuCW0HOfJfKIr4/k9xhdGSj5MprEhTsg1JPCDHYXWO5UbFADUwehoa2DJnN4c/LKfw6Lf
1nLMxyTN5MptYLYioEhkF9SSOh319MVWULZHIycSM4+LgDXfqOqNhfvNUqG2DUTe270iImHqs1le
bBn0viq6OTOsStUrdq50AOQsJRG6CNfpyfFLM7E1JC3DcTsPO0hwK8FVnpxjhfJnTVH7FhpDm3CY
LPBlAF+rM1wfG2KMfWSI9t3MxBIBLdVLsiZwF08gl76UoFxcCgqTtOt/797+pZvh2eAnUejITMPv
iDfJA85eLQybq6mQqfGFIuFSowLdtYhcpAjDHPJA0uEdc+Nec+XY/7u/7QCkgRszZTKfqvkgrJsd
zdwrXc6A0gBp4CqXnb8+jFv8g+W4UfwRvSur0MLeSUSr1k32AejBvZFeepH5WbxL47CK9wrZbCLu
ajLPygBPdQvfeEkjXGaMRErbP0bxMLNEI5dsqbREfa2u9OLbVEpHGfP5KnN9dosaF4/LRsvrSHsR
aNvh5KtiQCNkwGEElHmcYulWEHYwz2wMSlC4rdzeAarxJNxiUjE+gdSY39kXuRVsD346gDpUZO3G
evlIcd/B/QcPMngIAOQFRrGQ1jPId8YHfme7Fmqn/IoC7PObEh5sZY1fdNBlWDzQL5sIyu7AIf0f
ZTYc+bZUSNtVI9HjFm38m5hnml5NEd3pBd/4/3YrRG621OPjeSStJy91b/IcLGh0VYHLtUT0L9lD
Rx/Xl5cTy49+wzwyWFohYlqPyru7sthKV+pB6S8cbnkqVV36ltwcduitIIAwLuvSnyxGnHe2lmSR
L0AS0Wc9msddqkV5xnznsNgyFOzK985Hszy7Qb1wIym5R/uzAk9DQs5tnyzFk6IiNLduWYQm0gka
P6pPPn+56BLtlZEPAmo8T1YbwTa9K20x5fa7jGg63Wph7e4DFfehr7T9QwqWZenRlX7aFgQ2E+sY
oT5qmh28+RvqFEq00ahJX1M6QKie/L/IFZVgOYuqg6IUzTryAAOsteGs/TThNiRvViNbtvp7iES3
0sfaQrw1V1tN9ZN/bpZS4UU2Ma8IjjHpYo2IRK/CzShLAbT+OX3hjPbsvfyMyn8QnbcyktkmKacF
0F1WvmTP4xoNx03AkHd5tjVt0v7c9ANnhEaoASDyB8PbQQL+xPaFBkqQm/VGu7tv+K9iM6BdE5lX
r8me6uY/T2VGsyTdfKZnJhDBJ+/JW6zoT6XkQZKzEDVmdrK7Za1fmO8Ek7tXW1tllBPjGSTmFOgp
lYNQXymHSQkN+qkYSzLaUvWVWJSeumb1QsKvUtJGZR8TQfKak8ocuvOAAuKmtLW2JY8SF56eFPxW
+Fme3s1IaGSRyPrXyvQSEPOMGvYMx5DqVB1ohof3UwFTFaa1OZUlBAmF0oR/oVZMv3EkTZyMagQl
iDgMVggpBaTZvWBoLRHoM9W9cAB6gA9lvg2j9i8ak4YBKloHgREAsBuhAbOWnVRtjjqCvmSSFVKu
unD4n5zvJIkuh4iXNh7topAxpupLZC4NEDHJyJzBAx1OVuBDma43fZDV3h9oXTb73Df4Y0s5hfUD
2QawepEjQvJ4PUgAucUkj6t+QO6t8rLDEYtnNyzEVCByxkuxr5PHs+ZURbaocP6vny9+tP8y+LcX
sD//qGIHQOZ5QvhAGH2lpgQ64EQuqxCwtW1Zp3bUWhXrp1HMD+MzLBQ7yQGe/5Ou+LHcHZ+Xm7nB
4J4jThFcxxiUqQ91OY8kwNfKiLl+uRqEnueQDErF3ZK98j9g6tvB+dnUq9k55Egqbetlz4eEnW2J
RH1MEy/B0iv2kU9gXYdrDg7Uy/r8JejcZqD1XKUF1Vu/hT8154JgbJfqWJRgusJPoWvnzFwv0INb
Wy8LRskDyfdbHCKKdi+OvLLbUtkl3exZLP6nN/DDOYbvKIQO7AWnXOlSwWqfFw0kSJ8tHSSBwUf8
/yrP2M5/yviyN4sH/Hpxj9QERytrpaw1oxHtU2r0XmPZVrfZYl5UjFmgKEUhWGD07v2QwvGbK9Wx
PdioYU1P7Iyh6oKctKR2qhJTcY1L0gybGTN2lNKWZHKDP3w/3Hlm+9sJRX1UVauMSrfcsGtODzSB
JdRL0opjFxZqlF2EvxtZogCyOAzEHA1A3Z99XwzUJgyMRK1WMIDTr4JLft/KDI47sWEZRs5flKTa
Y8l+j0YU5KFAi0I+chqXSxdZvNnH7WXrB1TZ3/E32qsYhqQjcXAM0zhITUEjfLSLbJF/etbMVFd7
YJmjgFnoEUQyV/7glaR0e027NTk2KXP3niplM6R4Y3bu8UMxZeSKvqnrRoxTAE6As34igcPNgsbP
9GPvNB8G5K41kQ9yo2gNYYHnDd406LqhKI51KWXSHORQVHWi65ksjdbqPW3B02B8zm2rOL3WVF3m
MPEH4ada/mlk4itG7m3wJ48Is72PL8GrgLZrl0I482Fp4ovdsbi4mMDup3rvkmQFH23eHPGkWLSa
UtlvR974vaQsOCxivv8PVgNyT+iA5cd4poIAXfbl7AvsMszEVYyupWuEMysUAm9rWibDNMHuL6+v
4FHb1PSrofol4w9KTnt847/HBb/IObrHKSevXUp+NUMQS14GVX5kfPCZunzmAjG5HavJr3S+R9mc
4M1693k/rCZQrEr73HF9zfcQqdP9R3ksub6WFxRlhj2/22qBl9mqvtAwh9N6SVshbtoLyYo2OZV8
BDcI4LPhf9QC4bkirQ317I9kAUKz1oHO0BUfL6eseNX0ysmrPTDlizN02KzWS0WeSt6+YZ78W4BT
JR9tguehOuZZr/VNYa6aNKG2X3+9sxrRtTcAZy1EUazO9SsDxf7oOpxdQK+kY41+V0eLhYQutqXu
Ww8sP2kqiwSs86OODDOy2FwBfKI9yarrIoqTLVg3co+gWRFFbkUEEYPqen5uD/qb1UwwQXTDJvSF
q7n/XsWTvepix7wTef0jw2DhL9lQZELAyFzp2t7K2ivhh3OWz1kDg2Sjp9uy8ZT2qpz/qbEyTT+q
h8wrid047XfHwkfG80ycbXn/of6Q0eIEh3NfsY8KV94YgR08hrgZCxbMk7r3LhdCtKAh/3+t8cUV
n4UqCHoJeaDHt0vumRI0ve51OuJev+j9nKpMHxwtrlWEf/K3kuWuhkwh8TSclCvGyiCg69HzSl9o
ynuLURwncsJzVpIV9fo6XLvRHFcPfTfkNYjsgbXVN941j12ugHsl6XfRn/TNVP5rdj/RvvflGWcY
a/8rbGfMw7RqpMGOcE9k8jY5GltEsqqPbfbz6kCFeiKCGXAv8YPlK+OGPVektPwX9N6Mnagfqyyt
2l1kc+SuDKmWWfc/Hus7eyHCvQk4Mt4CtitoIkgSJDm5WYj1jqf0aD8XUEq9RVQ1ZdSHSmmhnn8R
bkYyJZy2Ud829l57sTwEGyJbSHQ9sHJeJpsjPCDZHvTGFZesdVlKZ1V9aSrZ7n4Jly+VJ9oGzlg+
rkGzg13x3BxlQuJyp5pLDxW7DyRIfZdMWIj4jlhpz1jKZs9NL0e8KebjrYa/HRhfyKbKcRzq5qKi
kbTSUPTOQZTJWk1f+Rdh9EGWwdOAk6A4DG2Z5qjnetVEB2TW7ksTmvbPCX/fVVYEhJuvqZJgj+/F
ACgRiX6MsKq+5fBzRBwkBWYs4tmiEolfm5/Gq8gB6EXSAq2ZPh+RL6fzuWcSdS+Wkanio9YC7F0F
sIDikgOkV9+45yT1m88XWqxqf57aZCXbDcg9+Xlf+BnxXPVrD6cno6vMzI+9KhmQC4WA0PtCjsOR
9KRC/+MO2h2SY4D/7fjY6BkkqweDlws/miFPuVTPJF+g9YItgMF+Z8GVk/RS+ZkoCrzV9JQHj/5C
OQOAfMCbegUWSwsUZ9FHlWrQlVNkFnLJPRBbLbLG2b0qqenwLt5z7kv3Z4GY6hWmL8cp3MBgDM59
xgsXjBWfzr0kNKnXt/lexnmc3sJhDsryi6M8kNdQSccP6dYiSDH5IwK7KYaM2sCKUE/bhEjlIeGl
fNC9DK74Pb3km6wFXUrXR8GsDfPn63hczhk6OAD+V6dXBZZqslKQiT4ib61nfMLr+d6YQnuQtMBF
JCg456EV9xB0qsQZeskeYWnNd0gT1ClrzUTYXU0v79jWdG3DTL+JvswlCj6xoNJIGx0UK5B6nrzp
TDhby+u0CDOutdW/PL5T0p1B/T7Aa8QBWueYSl4E4zZwa1wH8z82olRIfNjMzVVPlsHoD5Shx2gd
/RaXUR/QugttI88z/ei6w/sbp35MsUVqplNneB3IQWCsVvuychMXT1AknkhU6yQwQB099OzLG/Qy
EeHMvBzVmYAD22RDrCaheuQ2cq4BR1FQOZGfZ/aoYw8qFCFnFlvq7UH0JnPqOYKZRiN2KC/uo7Vo
1aaTJm9AkxuAXqI62sYZdWjkwMaC00DC2DCofxCYchw0P2h8blkNCvSODBpziZo2wTsTeZ5+E8Th
B7mvwRea6OgvTEoIqgDvAOG/tweQt4dTG6t7tknlZh/K+Xztv89Lb8cPBtL4ECoO0da2W53avKle
w8mWwzzpUkthWtaYrt/NtimfD6ypGwv4+Pp6CgfBvuYzqyRObMkyh3NEZ511ezVHxJj1viHq7kHC
Op0S8USbrj0+MsUmY5R2DtgeD+5KUFM8GirdM/Ie+3kMe8EC2kFk8o6XexLqjog3jevWPoWfMP7v
zIeRnQXF/icnkfcb4j3ipGbyoMoTyYA6Mvshcz5KXuRkAFZmbnG2FhgdgCiCQf0ztwvxnYfYRsvS
sqQObuJNHaz/cx20c7P21T0lzlamyvEBPGyXPmB7goF5blGB8nKQyaYuZHjEuHvhjHAAkY1dBoPL
rtEy2S86V6tThRXAYW4rtf3SusfS41tTbKN8G/3NFkIjciSY8DR6nsIbX/JFSDIIBVHRGP3BNuAG
J6CYRNxLWBjky2rEu5565Hq2zwAwYM8O80p7Ry88TEXnW9htKaeR08yxvBtERrooPi7N1n3u3Nux
hNjsZcpp/6YjqvqcOj4OZafrhnua3tNLX5lm5LCfHZ+YkVwfplUFw+4bWW2BVGldEc8I3aptGT8Y
9Ms763Nf4zB4se/obyvcuBD8xXeATQiUEEJ871yOqM+t3MsZPaBllF9MD/2QQn44nshihnfC6l31
C2vzhVAoXlYaYU8WAXo4ToVn2hI971BRYxH6PKuqJyLLePpsdH/6WDUabpXEOk0dVczNg6wQVfjg
7F6NCd9YaUstpAD3dZiaXex/Ye74nbYe0i7kzDW19Yo9VM9sy3fDVkxt+gdPUqYf5ucuZHKewWTL
7Jzoln6cMtSwHRLmTX4PnhA3ks7qnAxi2gx7bexCyYwM+UBxR5nD4tweouwN9uK2usKgfJv2tLR2
lNug+KEgTQvqvlP0C9rdiFdquhqmtX28Z0GZCxVSO6p6KyrQnpOYxUqXGO1EgnO8//eg+DgCvaH0
P4l02/ZEWXB92ccBUoSWI2lFDx6x0uCCzuSO11M9REqnEzLlcmySPJcOu5YVMROYobZBCErslsM7
KEQIhLW9oaMynH++IaVjiVQxPyWuBkvBtOkhwuhdw9c/zRfz02eujxxkojYShiAA4/oyNqBzXt3Y
GYJ8BQSGP3a5OK0MdTcLr4gQsQm6UpvRcfoVS7Av2cgqjslMXBAnf2a2qNk3j2GPAmjOaVOV1bQY
8Rg8wXs83XXcFCjxtoXejoISXD5PsNaeJdSuGharsOm8DPKLOxV1gei+kXanSrrCF5kJXdCqvqXO
cPm3cHc/QPGN88LzReVtMEy8D4NbCRXl2MIj2WnlW+IcigwDwfqhjCtjrQJsDNc/OTVFwNqe1dVy
TyAfElIIzgRqY0LSu9vhDcEau6ZGZAh8FdBfpliR5H5NhqeB6RBt9wnKXl3IibtuCLcPMuKLxY4N
HAceG63bH7GwO9oJ8pbLb4/jF3jpgir8pIwKFv4fKzB4qEe+hSpTq+VTik2MwXKVHIhf3S6jyinx
2xikZ2Ia2RtPxMRyDZ0HALUES8V5aL1ZqCaC6ZCpaH0IQPHGlAgh3k5ojlNeQYe50G+H/w8us49m
P7LxUsmhGgqD0yf3FGzzrqCHGm/huBAbw3M5FdLPkTz9ASvVnX3y+FCp17G2aVZ0BcKsMlc/pUPU
LxGvRNDAZa6W8/TXbAZNec5vK43Ot3pYPmmASsi4w3lMAYYunbWDt3dXvAetopeDery3rVAvE60x
8qhx9nG7liASWXlwQ0I/Rv9PnK1K2fvQdWgxQ7yuqVByAHvA1Pn0cOJG8vap/QIrSwgf6oEue0p/
gLM/bGcZUHx+d0tCE4AnWQuGsup6Kgrn2V/Uwkv7y9eMSJFxOhINeuRcncrMOOO2gx9yx4407zDk
eSU9RiHw95Ey/v9YhNz7AfuFMC8rX6maZyygMZmAgk+Zs+qRX8Hwq1vv/SDX6uhYPrRb0UKB0xKM
zP80c/cWwiNkvnnfnpbU/sC4l1SeoUnmhtctDNWI4OYCUp7ymAr6gaXYbTunfH0oSB70mZ1+sPCA
OWrgkU30MdxMcMPWvmZxuCQVCVGyic6gnksfKwzgkJ8zjrq6wFWRvQfDi/iTZyphR3pNFjGP8JA/
wI1EN2uVoCDKjxqyVqke92kr4PgYMasAcaGpaVNZ1UDQmVB9BLY2yakUFLWCkenDanQVixEGQeFq
BARcPzh5kqm0JidSmbaZ8Kh5dmfHyuxBKSVjV1kPGs28oeoVIfo3DtJwoJh8meCLOEJJ2iWpIR1L
rw6kp5KPjMmcR6eNQypiGbO+w9CoamrracIOBz5wBHoXIOpf5NQB4YFF0z/bjcf8fmqh4I9DihOg
zirODGnkfKkJ0TAkhioCaSYh9APpEzRlqvPfgAng00IiAMLQcdN2c45SFmIWmOQBYGrv6qCGo5z2
8OlXaOKGacRjgiMXxXw5mw0L0o2tQ26TIJKw0wedRQ2g1CFcXzi988jtgnm9XwHj2KuBncRE5d9n
eSvhX7coYI8InqJte7Ri2/XmgOZzZM7gse+aCl5UYuN9q5WtDfTv71jnYdM9wYWSYpNjyWGPZUDQ
PIk79qjtO76NtfIHakP1fo+napA4lPM1ZVDcUY1oec0y67shhTDmZWx4pYbyczil4x/q87ryG21x
hqQK/vnzQKa8HPC5OGTVFFRxjtqQRWI6zYdo3KJEQ5rtqE63MCGTiT8CtK2iUEch2kUwgvnUjrDO
64qB0oHjbJYeFu18QMXmWWqrOKXGz+YCspYK9gvaYPcxVCciF/UzBxNvo+yDPzZG1gA6EQmOjLj9
eSuYXuwtO6Oq1UWCIWLNtuyIsw1JhrUWQsA/9EYiq+ZDv5LNi7Nl4ugi8v0W/PFi86MUzp2XFKrM
YRQ9y2l14L4JCP1l8Ry8A551QCGXRcIGskTa8BKhuBlWi5a+CMG/3JWH5cDdU0uAGHQeT3ILn2u+
IGi6Yy/vhNUy+up/fRwyuAimhEZ9pbhuVl+o6Rtq5FzQ+3aXPyiomXo+3tqDvxq08doCt/1BX3l9
J1ySINnCPB1WaJXB0tL7w2dVSUbWza38qMRVJvvel3TEeeeC8kW1lEaIhiFv6iKdq0fIfv9oTNQB
toUizEIK2ht5setvvpoidvYAPIZRnmFO39VBtn0QpwhvsW62yhOEdWkkYXSzwu3gcdo566MEGhty
3ZuIOrw2xTEhdvjJ2tMan/fRG1oFqq+gBNB4WC1GPQzQSOY1pvH7/IsjeNS+Exh8Tyquxaw+QTrN
Wmqtk0IZLP9cJbMzVZbxwm4qoiqFga7/VAJSZBKAWm6U/NFxNDJ8l948q+yRkPKVBdoNr/YsRmSv
rfSBeRSNx1KkSOYwGTJtBBXNGgyHYsWWo6lntaVCd7tfdMjrPeW1vovb3XCYaVRRCbKpeOmrER6v
rHkWQO/K9xqCxnM0CQcR8ls+qLJDvd2PDAPzvaTlVD6nz/gY4bpiOC1lzgb7Ajf7vzrrDyGoZqmk
ULMrIFvjG1IKtBMsZRs5U09w8sABXLLqzx2Wsqmsz5NU339Eo1SnBW7AvojRtX76HdXum22aek6J
poK4BOzqaoEVE5Cz79VGiKq/nGR6+kpTL5l6b7yufMButhqILapmEm5H41xhLFxKBLnk39w+ZrE4
nd/5UOYmqAvBpsnCXBML9tL4wncDh7lYPHnzOhugM8T7zj2+nDn/mrxNSZM1hd5vAfgyZsklFTyZ
3pu11FABbk65ZwAWD1J0u4xS55liT9ruyEkp1POpR2mpvyS3IXlCo+LHIPcsLfB7mkiZhM9YrFiD
m2jq8yeKOeNQGq+CMiiGNuK1cxlPGm0oV0lkd4hl8Nlj3Wqx0S7CZcVRgIZ2Zc1G8kM+oYBb/ZKg
0SRfsn7mPFjcRDH6c49hocnROv7oWIevNtZFwAuvneIsEpK0OJAK3g9SI6EHJkaKaZhG9AayzmFD
fcaBbyHDD0O5IdX8Al2Irg7vq1kgCgK/7/AraxsrF1zum1WEMxUwRJ4HLewU8rif72OXDGBf0ZPw
sE02UDMOsv5jiXUrHUnSkee8YIrgS4DaOkKVr902eRB90/6HCcP01YLUIMvtekmHbG83xeBtgX8x
sEZdKdnb9y82hdE6yHCevFg/psZI2KCacg8YVVfbE2wHhEKIUHSfpNy+YFFvjJRL8AfULOO/1LoJ
oXleHaUn+OmYxybXAJDQq1pNVkqG2s/GEPddl7jaYw/WIrTmsXgjqCJMjFznTcMpivD3JV0IcHy9
EeD0LPEFAdfayBDoAvuWBVf1bkMnQGkMgIMirZxZd7gITTmSbJJ+1NdLV5BNA11ehIpVeoNum3DV
ctHFh7EinDtwFIhGn1FVfux+QmThqeGwkjfrFJhnvmYDU7RdR6xh2Yhx2yy24BhSN8S1LZIjod69
Em64uoDVSlso/HPaXCmCGucfHFOpFpozdgAcEJWD8VOxDjVS59Vk5ICrjlo2DXu/f19L4O0oYPaj
3gyuy9C6od0rdlhrAxw/QLtokXtq3OF9og2AzB64Kpz9IeywKe3WFhuvdXX17r/xz243fobGkDZ/
iopVlopl3Radj9k2lYcyxW0LI+/mZjJC6DzwWGE8fp2X65i8hrbuEH8eMO5DxZm1WwFQj+1FeTCl
+t0Q8I40OyBDFXt1zmhwdRdEPh9SgfoM5DydKOcSQIl4Fobs5D/crkqWLvX7RHrL5NT3sM1SR17+
QdJ3HvNs7gBnjDPjsSlP5mgkRlJPaAsyXw2/IcS9RBMDLm9jsGENj2e3KD+Uei7H8qLFefuSm5H2
DsjfwX0+hmK7gZaRpcDNtafAQIiN2fH3JOsF5mzdxoTdAEN8rHxr689g/WpSjH6rPIKEYli1Iz+t
tsvVOlYiSAYiHSRzhwFUUAeBjSqs931Vm7pi0AKep+RzinzEMdxbViRz65nXx/SfUVkYtyWaijO3
rAsHEtXJn/S5Kao3hbUTKPvUlRtR8W/mdaa2mHG9nGCuzQiR6ybZBKJuYqc6W4oF4FQCLB8d2InH
vbZ33II9dRVI0+cZd2bwkuz6Y6KHi0n+sgXgMfK2YRRn1f2tQ8n6tIZd/JGzLLBbYHWZUh+MYK2d
PUz7JYNYK/BnMGHhbXjcLWv5wuU542OTB72SR+HmHSbIA29fJhoz/wr/9S/Xll7jmLeDDlwHnpJi
Vm6BPirc8UwpquO1+ihRcjnpt5Su9OpivNe168RfFuWYg39ErkKZxoTrh8Sf3c95WxOgUzEGfhi1
nZZc8nljTdPLAV0RONm4tE7znsl17a8ZXRIKbx7Arbs1xXk6BP7UDsJJY1qm32oVQ5mFUI8foKBL
6wEAfeKqL8Mvr0jx3bboomzw36lMsA9n2rfiOvvk0I/tnspHhPM2gsJ8+JX78SxK/TpnlvJimbpw
NqPAXA7klwHSXan8ohnuIWtBDVd9cGwY4SiDKsPepEtP34u9Kd32b7y7MJXi8D3Q3vxVg2+UgtDX
cPoMdNAQCAgTR+nIUGROOastAgmuP2UozrQW+ecTBI7y1sSNzzIBK6pt0IxgKzROHpIYgy2EwAkN
mNReuQYchwwy+JaXghcrkhwobRwqabN2lP3WnV451r65xEbbSh9/o2vmZelJ7AFVBlvHG3fsVgaS
vbMmIhnv1lLmoQGk+jKEDCCM2tZBF/UpCaBM6Vo8N/yzl2XQYcpqIaylMEokuFuCIgF0U43L84/f
TojJLBaB9DXKDv80pxIBDQmLLe3UvfZ3Mu7D3Z+pfQDXJ/2xULnQdOuips0KOCdxmnRG+if7SZmz
0KJFbP/uOcqTvCySis7uJqZFa4kxJfvWuOc3z6Sql3XayhFkuk6N8UFYo76sX5F5POMSnIZr6zYu
8q1wW4Llb6sTxCLHtNvHrJeCviaOE5RiXm+yzNb6mX02+eBDFB5ULREad/BHaz2qXm09Lz+7zrLb
NOo+RFnuNuUAKfWJERAAnFcuQf4h7+D/yVJLpnMYe6PabTozx2KV8zip4JjQPjqDR+zDqZzWmJ5a
K3mb2WHCEtXGTYsUH8wwhtJu+jCnv3hCVPXUyzsEs92Lu+a7ypGQfZ9NK38DxIXOXZNzHha3mjJq
PbLcp9I94U3zfjtcvGi50AY7JFqpecne0I+4xx39avJVu9A2ImNX+9AL2W5UkqnvZAMqVxMPn04n
2jN3YO9Agc3QMrJ9wheKmf8J0Bl4qGA0QXbqxJ0lNv1IbGlrecBeXoby5ZAc3szDyUp0/7yZJ8df
sho2dRTBmMctzAkOt2QIKGsWQ+gHvtbtWUTnQY1irA2D/X2DON7CPd9PgGVgc2O67e3S5jhgYte0
uEQOKAfnTBztOE5gEfi/PXbBmTBdNdPC0wG8vDGeOmpWUR8B+FA1Q/MnT+qtFqh18ll4RLeY54aP
mJdhidOU3niri+WQpmw1I4RsgbAK8QqBjRqTkfa1hfxDAVialMaGhm3U63WWCGX+O9LDIWgBXNUR
01il56Eus/BaTqrTmYqzBLU2myyotL+04jGDOxwJoS/XCp7IHdYKPMR59h54DRqd6Uw9a3mm1P6h
BTsAm6VYL+ohCXvAFB/VSTt0X5EcoE+Jo0xgvSNyyuj/2ry5Hb0QUjVb4+7iTtegg2TrnU4kFazH
tX3FV9EgDlGRe5WdV9wJJ2bffH7OAHHdnh8cyMLqkCVTjtp8OGU5nQmilm24dc3z+GduSLwt5DBC
b2I2/L2PosReeiFI9f25oMkYpWaodzGrMwpsvYcQgjQUNjWXhJAcjDpo0ALeWbdhMhwy0FN9PtO3
AyZGz0R6lcBTsAO9XQ7dRri/VQRpKP04Eh0fnbs6EvGEZ/wIl2kWcZcIhvaQLHPlogwQ0lugm5Xw
kpvYSr3df7h6gfNv2beuiuN+qEQdZ8wZt2JkNN5+PdV4gWSq8EABFmJ3ae9evQPlu7YS4RJ8Nv4S
ErU8ynEG0EadCA4pHIc5tHO+5w36zwiZE476sRu0Co/gq7KlJt6crw/wZl+lzTGPYTTlH3J1Hpki
F9v0Keghf0xO2lH4Mc0J6FhVO/+Cb1W1+UTXUviL0AUzQ7laOuoxll5Q7E451mp7MC2uxvZDUna1
sAR22Zg9q2qF3Zh/nGwj9QAeBt+UXevI9Jgt/8FYCeEfL6bRQXT8rh57Ivj63iNfxNISyMFGpAx1
gnNwFqdLoMqyvLqOG+U/8Hl0EpJKeJFUMKt/EwxLmS3cQT0r8qt3UJRqTckHo58esvjdVUy1TwZe
JxbfWhYMLMBNIceQ9bCRxaX+MjBLVZP9oBWyHCGNHzZnHPVYG8lqZ47f5vCwTLCXIegeBS6tJuyR
M/cxvR0mtdhkTqIcbrJbknI1hCMYyBTD4A1Ikpb5H5gA+Y+n8D1SJoKClYHSUn5fUj6yHoJkZS3A
pYeY4i5cd3Bgugm1NcLhTjD+//MeiXly87m8Z6mIV0VO/aI1Bir1+zhvqpbfN8VC+k97e3pd+e4T
ZL0cLb8lCMTZSPvBEkd5rwBVO4e+/BmsEnmL80IlB0MsdagGhjCQJ0YikUmSctSV9AZI/mBaBzPu
YNEbyB5Vv5F/R/uYs62XX0ygC9O++83A/FcEhzWI62y6ZGgbZ+bok+YhE0Lr7n5JVhKNf99pnXFK
6tVYJK0wNZmvOiLnkoB14a9zHp/w5y1RCqQ/qMgDN6AySJQvk7T38POmr73tv95HzuVSaRZnygfH
6tS686ZO/dL1MjaPwnYcw/cizjXUo1TNzDJ927Z5qaL3IoYO/G+mEhqPpVukNR7KUUq7t0mw+zLy
keUi8nk05DVBSTcPBrDaXmyVWMkceupTS+kko6620JET2jIo21e2WItxVN7DZyX25j3SyJfYamie
OTaB0zvvJVMvuaiYH3zkx175660P3uVBUC0SJWqooE61UWmRZ+vRxQly6c9pnI12BxUFewzp6tdd
RHaOBonnpAzO4yG5p0u/5xp2FLF9gzb+MK6zHxyE3TPhJlzeiMdKrafxo4mxRlvlANVLA6iiRXPc
bL4ff98wiz2XSIjnB992IELjPuAX0iq937ulmQDCkYL9zmRNW3NrxdUdXquTcN6wIq9Ok1ZgC+FG
qJg8EhlNTCXxwg6/hkarNBPlZTopygU9DCCIc7ONIBHZMxJiCc9Zl2hHSe6Rp/ZBSX8tLDQ0Fbt1
DFgB3ytNgdp2KCYVn5SyX6aevQe45GEymQDc//UH75HyaxS3PrfVtHmZy3X4fNnmQ5gU2UnWSGAy
uJEdreyET+irsi12gGv8wPgOHaTWSJ2D78MGN80P5lORH7y+YL6I48k6WWCpDlGFbQ0NiaqFmoe7
aAht2vzSmly/gfuRGQRmcfFFKD2Qhs30oDpe8zfAf3yi0zNyn/nIpUFCmYhCA2mIPkRhtK+OBtP4
kN39+NEvw49ZoMq8Fm6zBZM1xP+fykzFtGaZl7bJ3ugUSskOMx4JQup/ndvblcfZbG7nyF28aGCH
f2m6XgheIui6O4g/2s/HFQOcZ2hrpUkL5shROUuDO6dhI8VwJJ9HYO/L4yEHxHiu1WcebPoIEVV/
e2NjneTeWzc9Pbr9GDqc68zBnl4IcrOZn842m/4CIpUTamKM6Xbw8I6d/LGVvd8YtqvD37mL1xUb
IuRdJv0aLOYHxZQkZVI0ekr2UUmKuDVo/zN1LuacGu/0LV/mIdvyYb2lC47qa5IkQgywVWVJWkN6
qxW0PY+ojcDG9reVV8WDSADodRIqKa1ZNNb1EYbGQIP3dZr9jvlPd3wSXObVMjmMQp+sg9brS/oU
hpI56x+mBviOH2WatUYurCV5wGpklLb7GgYI1a15c1T9U+Kmm0n3BTQsXOIa5r/D2L5dmlGr33AH
Y4eAJHeroJHixSiM6zUgil0utNVR41kJfMHxmM/CF6T6VPPziIETpHvV3wn1wCVlA1CR7muovpsW
KG14+l8QvjYdEu2sw28oX0pfbTgYpR52q+iwU4+yZE7XIErqi4svh3JiOh+N9t0KjQSP/j8Vwuad
aaVWv7LAguiTZw57sajiyIt5/gf6OxxT19J+YSN/eLIqvU+i33kDLiI1O3IvIIsKN+wQXqW/Fu23
oBQha+ymvvGQ5A6DM2PqcDDnj0bVSKsRlgB4MgoyIpoWkKJxX7puF4Y6/G+KgEkq61aE+6qEpSb7
JcN/Drd6FbmHCNJmVqqZ2ffqu69t9rCZF+M++Ctn/LAinB9CnEigfajRpFLt9Ev7HTYdk+TDVjbZ
9itZ8fMIk9rfbWc8FqefLluyQHebApJTv1w2SRaz5kL3VffLh+g38L7xqzSwNCSibkk5bZl2qorS
SLB5jHQ0+FbEmGRF6DCHctM7wsl2TasWxbWpYagbGHgis3kYbij7Uq7vlPct9UxURDQfqYMiuDqf
gWd/dSe8gu2+o1xII9OBzXTAr0ulryUMLQiKuXTkTJGUG+SYoFGsYavyUN3uYF6mayhAWJdQHfcb
YdHivpvb6WHiN36fMbiGzHdbdOREhf0FO44pYJQhQgyFKu44BxxOS36l22SF1wh8lDC4YvGcLgQQ
NT79rFK3I3k+34SumBZfs8ajqCbS9AdvpFFuK4dpnT2iO+Jq+i006gjYHWsVHMzB0sM+SdoRjIPR
dPxZTXRZk/8Ij6zmRfj7yuroyqcRvNKXv9RWdrCNthZ6poephE2FcGQc8C8T1h5n8B9VhfYtn0Yn
pcolXQbpygs3UqXit7O3gsV3gIx8heFaR/0DTxb6K4mRI8ITFQL3N8rLFV5UtA9ivPcN4h6Oc7d1
74P3OpRDkCBYZR9Pu1sPdn5PmKlFRQi65kOpXVEiYf0UULBmglZofPrCqhd7LN0zRG/Pq2uLVfxE
zk+Whdhl0Is8CDsdAoZlBMnarPp7+LZ5A1MRPEOc2bjT05V8RtByztHZORLmmPJpEDRf8h3C+w5m
2dAX6EhpVfygtyr9APQ/BxDbKIl0Nv7r+ZVtZlaE+gExD6xoA5YLEPvZYWLcNUtvQonYJqJyPlea
aPwqiLEu0vHZENb0uxonm4LNkHPrHUzpBZAdqAAtV5f+tD3IygAhtIwrcfgzprNskwH/qwCoeJaE
wCoTKi12GY3hMTEa+t12qSw385QJkIrlTebfLOLXQcQlQ+YGhrNl+bGthB7ll1vLtQE7t927GTQg
AJKo0TifMCSqFde4wJb/9nT2pgXfs2f9pHMImR9HvHIovgqJszCNOgYyHBCrnMux3RjPT1p86mzO
4G7Js/hR2JF1dmOncDMHIteoYR5HDoHZFx+nHxixKn7tYClWHILEo70Y/sGIjDXJzkDZLEfLRrMo
i81gQtrH5qK6gFeOxi0oplj6C5lfVNIPQ/E/lQ4/3z6cjWaZp5sgcMSZrPNbDaETo8S+/NP77EQu
Jyae8KYjmNJOl5l0DUQLhB8JxdDbwp07iScLiYncVL2h5LKtbjOjvFBTKBVOwuDBYr3/Hu3MxQPR
WqfcOHfC1S+r7ajUi55Agtf/VcaWm6lN+s9muX3Q1L4lHbuk+iEf9cKZE5BWlna4n9tCSxdzbN2O
LjUKoZUiv+MYF3VE9wtz5YuTtGe1y46juiPvWKx8FOLDWs4ZlESMkKfj8dgBXFE2RM69EsxvTx6e
/GB1NBR3jc1bGuJiCxVlUvIdSL+flimJ6nG3e3DZypa61dfwDPRLRworfNfAl75x/VhvtBfGfdzA
V5vsSn4YoOvVg6ffx9tWyWB9pKWLP6wTLI/dS9adKCel7LLa3nWYqkrISC2x+UcocCzFA4BXLrpb
kCqu/zPzv9w4lepg9aXIGOIYjuxBHfpkHswLZa/ft8gEHvDSKtq184WqNrSLI+oVF6I4hqUfaDHo
2sk50JvOLLguclS4SEe6DgjXiv7n6+Et4IbZiFbPirBld3R110UTI/x8vpf1+zxzOAJpVxFjaeFD
VT26/7fI7V1EVMz57hWX62M/V60tyTiiiCxfPevvwXmVDMs/30WNruyGNECUV+OIhwl8JP7y2ULS
KuOzP8ANfdntYjfPyxfG/wowxjHRHx9wBoI4f4n/WEsTSg50jmuWq4PLAtbPyXvDctf3n44hdJex
T8qTZE7XNMLnVQgcATyhi/7MZ1XUwyakIfIeGVjXNw0QbVno4HC5j8xgMTjwqnk8Kb5BIac6RTQo
pZJMlLWgH+HbdHZFTESEqeZnZ79z8GVubjHKmLvHpmCt9HKWme1hIfdsGdXrE3wvAI54iOTUbbwz
a3bbC2WwJx6g+WK8BMhlfnXqyBu3bZOHolPxDxoJcKwiPaAOYMzTdWa5IXuoM35EyUtl9H5HrApF
sb2i8X4TVJJqwXLxWH6n5fPYbZj2+4cKUUhRpzKttrD2JVWibWGCn7Nrgz2hNH/A4y/8nOOE+wLl
MDze8EdYjSzu1CKSR+FeOQ/cyjWgcsXK6I2YvLCTrbLGvfuHyk/nywWyc5/lsVEJu2J9tSBxlWA1
zVj85bzykxhiWZKPoU9GowI+FD03pXy6X/QDwXY3OAMAMCK/2GKtUluBLkyUOn4QF2HsE0QBa8k+
mfloT+ut0oHqXjgbmTGCwEz6HJdCumYWZFDY0uzR7rTblx7IgCONsw2SKyduVqYpUune0FM0SoVi
58bYfTcoebmXx0DyNO133eoqknviaJ7kjAH0/6Ao4fPXJ5qcauCL4Red3wEkTzCSE67AuEeIU0yX
fc1w19w24oWU7olR/vUiryPqEv4clB0zlLp/ldSaUileg/9NrjD7nJwq/9ZXf45g9loYAlMRBhwJ
wFYLKfP2ewR+mUjzmiGGRVo0unY5dyV01Pp6wbRjsfZa7Yy9XiDFMJ4Cl77VY5nrl2TrjG6L+J7V
nGtuObh33v2RrK4w7YdYZm0QRr7kxxmZK+u2nBoPjNo+iewS/749wy9/wdY1lfTe1obE0YV8UJcj
zDH8n3zmSa2cq0FxU8La2C0SEI1w7O9j7kZD9AckGp1IhXAnA2aeSfdeK/m7ZAk6eFExRlWI5VAj
MkhAr7Leu8zTubfxxo/I2iSEfrUoUVkjIlOqUOfveS6/YjRIwlwj5JFcgICVGqgCtW367izspfpt
8Y2wyb1Nu9Rq75PQt4BjFmiZTG1hlBKiPJSDUUHiJdKm8iz02kV/V77ZIBf1obPox3+FwzkEY86Z
5iNWuJSn9yiO+kh8vVWG0oOABNsii9DNM5He0XSGZxoyqBbYGwjrURtgrqP18uuITNQV3nZ6Pp/Q
IIyj2SygE+aoxk08ul6W5mrrW0Apo8MOcX93a+o95Oo0QwhD8L0RVIMwUZpY3GTgGG0l/EXj5hgs
maBm806jUtC+e7b9sG8v5A9ekuwyNgYwn8YgF0cFbE1jvfnr2y4VgJ+IPvMG5zgOQ5M+0Li3f2R/
NmkyL7vVh0ilOteDnbFbyJOQS0XXW0o+wL6aqhGcC1rMPWiVWkENqqe+xTrVMWD8GtAYrEejtsRl
ZIC0Oxueq+rzSteIlZOhxSfbHadbwvDFIYSREaX6vKLwrC5ZUpVbHTQ+nuPXU+F9YjLx/usvrXP6
A/T2ln2OG6csmX1nxWogrq4wQulZbC0rq9sQ0xe2+y1u4OW1qjlD3e2wV2tLXK6ovHZCB56HIZn+
kwx/iu2ekZk8v1wIFNvCakE9k7B3Gsq6TnCTQEnOI+kVAooJvO1UPYbKfyYlTXNXVV8E2E62AS0b
LhLx3yn3eohTnqxNEITmQV0RzIbUgjEZtQSUEVC7NFWZBhPTsnrx0bkC5cTNZtIbeLuxlnFBj8kk
fMJjwqC7u5sKsiFjkTYQjPaZTDY8VaucA931EGhkrlBgIONPqLfDsWyvGVoFnpYp46l8PF8vxj/5
jS5NbRNWz+ILXXN/BtJbTprkOMt0PXVneQCz7vNmdX5jo/VNIt1/UqoXBTD2gFD2XY1wrbeCAHRK
/q9DaLVx4hf2ow5BfB7UZU6TIs/VAaSdXvFISM6zY00JNHVPjtU/nzTt2MBu0KW7kzVe1UKYAKFK
AwdE8m1LVeWOLarwJ0R3u/io3IDhM+3rUmp+iwWXP7dkaWa6IuKvssCgZHPNO9I0sCIrEWHbFBjN
MPV9Hs82QksF/DaxShlWSJOGI48iigAbmQ+2yakltxPE4Ay/f0LoPKVRnUYJDIqOJjJbnwMjZh/J
wzOKkFWtCVkBrQgDCu2mFzIZlbY0Jb49RqlzUxVZNz8EB5rwtDGIvXtFaYwHLceeQT50Cc4oMI0l
F1CNWBzyjs9XcNlUCqNIxRXodQye/MbMr6oYZNMS81tGvy8mLrrTx7ELl5OLirLZMTfBLOIgQDhS
tzuNnXFNREgKOndT/CW+8Oitqi1WJgjkYT+GzU71JZWhMLwTyqpJFhWmJu6oN1dEOeYRn557xJOs
Bd8/YjDyP0bMdj1DNSAMzcxmrgIR338NWcWnBPjrsHJsGjazFlflhrvIgk0+rkNGvvZXJFVclaR+
bNDS6l2JML3IILlQ9+K5fdEplNZ3n7isvB6JxjmQCwcevgok55IvcUxGNQV0dBNMpDPIriwMRWyq
5bRB/HzwhcGQXtWDfGx1WUtCcQcG8KmzBe15UCzdaeXt9Xtxv7L+6Rd9n3PmysfS2jjLDQcGn4DB
fXXv8nMb6XSYxNfxJgXGLiCZAXPGXk7I7gTxV0ad7ssI6jlHMEuPSgC/OH/DzZSYBkW0RJKKFQhK
4jELDMlh4w2p4vMX8BtnPYFmupzNnogFZ86r4pIZ1SfQu21q80coJzSOH8XyLSKv6ravL4JOllOS
qJc9J9LgJZqYQ5h6kFb5L9vZ12zW+8m457eZROLwC0uD61cLehbNqxHXvKzW6a5vXv2lJNsnsOs2
n+vwSvQktsr+Rp5of+wPrarYqIR4gDHbi0kWFj22OJO2BaogVF+vnE7rwFTmeqfep2i4LlgNdN+u
tQS10jw1KeBdwt5a5kXt1p9oWWRmOovMe6G2QosJ4xNFMwnAY0t1pO0/3opjOyW+dejhyz/pekVV
croqvYaTtesHLHiseUfem3h6KFrykPxOYGy7ZWTtRZMEa8bg60kyWBCWNPo4PdQqzh1cX2VaUq7i
Dmn5RwnYL7tBCyEFYLm/eDyyenQjeWWeD1wXWvzHhS1j9ShuM+8flywNpqbCRUoEqlEiAdFZQbe+
9AjLlHvIGQ3irBAJ23QVO9xUGofZIaF24araz46o8lrcamIQ1Yh2bRQlXPemnJiL8QLtD+fWkzn+
rNIN2Yf198f8uUZozv8rL7LSywugBooa84PNCaIY+xo9sXxkU99wbUZBgu8xUw3YePeu5Hgl1R7Y
8daGtgcgn0Icqssb543W6DRieklJoTV3szRry/7oKfic3KB+Npt9TqSkxV6oEpf03HXO4O8QROOg
n76Wt/gE3fH0g9CDADSXK0Oxh75ObGF/ThtRAC3dP8EGDuykMlGahD+qU57o4Wk8gxnWVYRRh+CX
bmIBQKSZDZmngPUlHkYfiwFJBQSpg3N0O3NYo/x2f6Rlhj7+QyPjAAkz03rI4sAYIMqE4lLJStKr
ScWJu2Htt+iUIDCb3PDqdzTuIum//3nxVfDQpjz6VRh7ojKwcu6G2FhgzKseRqMszq3NkwLAtVI9
jWb4yWf28fRQQffDbIiUf3prNiKi+wVU4QbTr37yIYrUOMgWk1vvXUkHaPy4AKtZptDLblgWkDUc
fwFqaGCH9AcTe5nMa36DOsVv8IrubGfUlsl2XtVJ5rL0c5JiCImDJfweVnHcUW/+cI6U+uwaQDmD
kYw+51FM2QorZ9RidMnknmALvdJusMP7TpU+ulfCgb9WjUcfPcsJlUIq49f3gKeUCCXCsVWKtfPX
tqkE743uQRjMh9unS7d9RkuNk5NNqjkVxMSkd3yoX/61ofDaGA+g1AMkZO59rsbqfsZP0u2w6zCb
vVhchVH7S7E6GNbx86TibIHWC/OVsclJGVdY9ZSnM86xkXXu4fxd4oDZqdrRgdyzMPhNYCl6bBd6
fQAumuD2MsWs2Y/SGkEDxA0GwtkkzOf2VR6c9TGsobM0uSjfl0AI8ydSHQMHDSUTbFH68ULpT0Sx
B7IQJdbWu/MVNwMX9T3vgQbQ2JVHdw9bAQbu2yPguQcVaGJujYPlPZtEofA6PZ6Mbmi+atgUcD9u
tbiOrg3OgPn4PjBC7HT1lvOMfgHVlj9kbSr89JF7tRwfbhXbr1UC/MAG4+1vmWLDoyS7ZczdMO+Q
Vnb2ahzrZt2fbJCL9emX75T9U2IfBJlxVbW8wH31bcdvjr7TB9pkXdOFSweyN8VF1D5xMoiMqbkZ
1JOCb4mXDNIPGViAYkrfJYo/uXuBcb/yNWUl48/Jtb9+B6MpMUOkGmsGe5tsPe1mndjuyhEpwlDx
6lV26lGeGqIvOwjd167Uj1O+84l9W2I8/FP/rnDd+nZG39ectHWBKaC/JTqUKDVdEDSmTj0NvZIk
y/GpxwcPkCGGYwZQgw+X6W1Mj+pKrNwGcAuTlAUmrkJf/gnLr9NHtsOYHg+g735dNQ1d59nyGZak
WzfheMfp6WzOU8rWa15muQPvhzymhDnwJC7DpcXCyB9G+TtsMr4Wdft44aYRmAZAuglqvjp7Ovxb
Cl2aNv424U+aTDl23bE05W6CjaJfWRMozjV7ASv+Jm2K6hRfgNAQbllBXnw52wv64jTqZBylV2FZ
s/uW416r0V+rbpVmriQM3AeIrJ4KVNAVlyJaReUIGChc7TgG4gX5uSsR0/0gI4DuHEMf/SN19qD7
y2PH59T7Pec44Obxq/7Ue5bSCQXI0HeKOO4Zy7FyoQ3JLUexJyEs5oSiiQ27p2vWAfo/XK130/47
pv057Ynf4hjGj1Et9u7bD8tfSWpcjZ09w8wUNXkL11tmeJzypsUAS0hEnHpoVq1J371tv+fTWyM0
oMz9ikOaBd2RYHrr9VJlQmqZ9rPrKFvqkOQ5azk/7kFT+19R2i1ILU5GwdWJ+UuSo0Kdtwe5HsAg
o/8/AuLcxzvexJ3ywCZHF0q1cQTbor8HGZul4JP2E9Z/BCCGIgCcyF5P+P5ntRDsWirREniofgWw
64+EwGygLBQwlf7WiytFB9bV1fFhumtbsbdus6/h2t8gHJ7cqQzitd9QENCO0korIL54iQcrkOza
coArks8hg1gvkVYtquRSrGfpyAsVT6ipheVug9HjQk3THIn+DHrov7/0TYAaCMbxfUdGWCYCTL6r
LZ5+VQ9bT+dsfMRrgD4rxz5KNeCb4MWOja9JYgkpbC4J/rf4gBo+HylqZVWy52rdARmaOC0OSRE9
7XS+6Ogyjy9UnK/wF/07L2CpGsvpjGs37JJvJpJvswTxEr2cAN/2ecwhv1VICIVrAsbxKZ0dmirj
QE1Cj1TsLSZWCi14UZNNeT636akjbMekOoVKkMoh3RsBMeXo+md5hM8mPUUnHJ7fFhVJNf5W8NRe
Xbx4wJ0Wlf18hbjGsmgkbrZj3OwpHpjWQmL1ba1hjVlM7B2TImyTcA/bBtSNkJL0kBFbSvum/kl6
pxrJAma45XntB9tLCAGOMoiAvVxQuI6ZuEsU8esgUt6t4WLvybiPRmW8RikPvXEzvbBMFnT+cDd7
ews4wYmHkkxsOXlvpTTopjsSFUx2CukVsjjcG2dpVaHkRiPGWtFbpjap7AUeq7er/NDbDI/Cm18g
ZcjzYhTvE65EPGM4BTxJKErfIqNXZmu4WZWJvX7sPt8+Ll0IDsIk8HKzZesTSuga+oFn0BYVo6o3
yPEJWKGXz5K2mDVODHmOL5OITy4v2qAJim0R8IElauWTvpSyJxSlZVBf/d/xy69dpSpYgcolcTBw
EO9ah2hekjGts48K/3+oZ+D0kRtYlwfeX6qbxv/Btkr5s8ZIQnn45bE2UxTd+WOaMulgaNse80h/
lwnJPCjvbabvX1wgrfaD1v6OjwQeTsvVu0b1wdeD1pbWlZaL/Xqtyw8u1XD3zQn+fKcMfDGCMrSL
TVRej34g7sPsUMrPPBsiJvodntdOTZGdBZ56d2ZITy1HaObc5aMADaJ3ImpNdZZGgetCmNp9xtP0
XUpThbcjU7D2CS+lSrmaE8EzLv8acAaVKpuVSexs49s8BlW9TX8WyLyZSnE51LI+PqL6pxkctfK5
E0uhejhulGDy1ALeSw7hfG3YLJ2t+w+fZhAlWtDMmjxte+igERRgIf6IniWfZW4j/BC+jgCRFDbu
E0Qb6ddp/lWrR8knk/OsdxmK7pg9T0uRn/Zv5Ww+E4XlW9uh5MkqkUHpQUdO8adqlRKxEU7vrD+K
suZT1lDeuvpo5wEWkNGJY7uL4Xa9C/gCAzNQlOv/Phq3XDbXUH8FbX6W6gqriJwFghTR1HONsMd2
hcqkEOpvxbJ/33r+OaAqv4279XgWOQw+fI/+JAypl3qTk6Vr5EuqgTmz5dlVgq/+WKszZ94jmZuv
ZvvzMmHeNV8okVw4uJfhEEzXXOYuT0msqOVtbLz2hm5vIitzFmoGI1xFDdojgvHarSMvW1mVKXhB
86thjvj99vb55+TzxVszGX+glXxWmuza3AaruiQq5VJ0BCUsGub4iJT86v25SC+ohZ5RGMOSStZU
lhBmfd4wF/Xe0qZ7x80ld4FmScG+Apl3/NWrjUcr0o/2JXYI2i2R7E6KRXunVfYfsdAGP2AKz2pA
xdhlJ3vC5gpiPvegvUxlcsR751HDuLHqZaqdIiJEkhWcyd/Ffa/kgSR1n+q1uTBkHx2iaaDmPoyC
R3AvgR7+rdv1AwBrB2znqutT61BPFH6CxdkOk+oerlz28sNaY2+SzzODw2Mih/1e4L2TCaOc8JB0
DWuEt7WwJQqGb72VtKUmuKpuZJ1FavFJuhk/HssLab9huXkeQFSPmHUBPAYBM9oyhp8pRXEcjBtf
L4EDx3MYf6HRbMdS9BLDo4h0eHIQe8wg47e1LDYVEfk2NccQXYyHItOZN+1FsohNn45tEwde8Pcx
a8kNFjgxLaSZkSUrCqNzksMjcK6wNMhJyjUKem2KZf5fOs70Wf3JCXnXuttuOMlcXBlCIhQsZKKM
YFqgKBb/Kpfif7sDeyU5dlCc0gg8YlhsDnioq+vuHi1c1NIsaiwmliVwF04tnxjDfwc3Amm9iSps
sOE2/vAyi/m45QLLAFBi1HrjgPhNUWRMaUECWzorFuw/x2kDTNZtzvlMb54N0qv8k2o6b+YB+D/e
DeVwtKgUFK/FLiDsEXhapFt0kEZIcJR3MnV/1bxnSjp0MwZXzYUOT6h9+bYrbZ5Uvqf9uf8iWsY3
qHvA2ydrFX4+Sqiz4f4LlH2bsyasAQY5PI8S1ahkd4lawJsIHKIL93wABr1qx8k2CYciS3qZr2fI
0R47Vlukx/+RE+YWU52ORrmgP9s8chDPUn+Ne43l+z5Nx7Wx+vi56JhzO0Kkl5Njv29Ig7vz9Mkg
EB2/kyP28gnD0Fgq3wxlw3ORYYcr3c+g1KyiDhLwadeRUTqf+1PHppdcWlVLOLyKgFnSn/ZdUFpz
hlhqVZTdcQLt5GtvkKvdwB+BTye1UoqN4410tik0Vs05Y/qv3ds7OAR71bRu7e/AeUKn+rWCRw5w
VbvicecX3b3ZXbwOPGLeQuf7jgPY6zV873dXVqz+wfmxw4yYjRDf3o/ZqGKFbiuGdWhyeHBn77Hs
KSDGqa/guUD0JA2Xryr2wR+V7c1z3sp1pVcSBUOr5djk/b6kz6oNYjA9a0YgUbhfrN2AGKWfXw0P
Xc823ts/yruaWg9fh7wj579NNW4GM9CcIPM/zRbu5CkhtUaxxkjieTpCsjCAMLLaUqGzQ19MBbaz
PNwEGD8GC7RHTgVvgaOWUIyw2vKOKHmf0iuz1JJfUAOykcgNLpWOP4sFjiIIgxrKjX2BxJZ7dnjT
PNVOPTklr4fIBZItbaxBeFH1T03mG/yAlB6yOMofqODvclvdikuCXCc/QeU3Cd6O42OASfPpAkaf
5noC6LHDqiP155Xg17V+JD784kuGXhqEMI+7tuQsGRsXKcwtsiwwtEHjENtE/+oYWtXF7vJuMWyb
5h1jJLzq8aQwWmQ3/w2NxMiXISBewA04Wv/N6Zs6nPJ1PVeF3wu9sM3ofRNIK+Q03Lvy9rB+AuG4
NVtR7F0CA4gSvcQosQ0q4zRg6CJNRDe4ypUsX3p/B7V3YcMhiRZyRlA80Qv7Y7T5ZmusiXCJUcIW
6FGAetDRcKX1tBzGBihyr/STCyg01jjvbTFp7bJ564pafZzGgHSlsyqEmgGkDbcF8vPSys2DH97U
L3QA7OLvx9gLo5r7tVsWuS2id3jxW7HCZNk72j2oQvEDxf9T1jXTELzzrDSjbkG1PHwjG9XDHZUo
0ERJSLUqd0la2VRsnaf5r43QMupCYHgGklAA8yaCC3xoLWHuq+W3aQSO5yQc3PXwuIhfxHi5za2n
6NgELO7l28rsxKesFk24qv4qK/ZUtSq13QhlPaWArMlzBls9U6P3uw9hasfMjnr9GzRTRMkwGRTx
94nfNIQPISX9WeOFbzntZdRr4IydAzMqzo1MBTOTUt47he6YLqg4ezeQyxiS2wCOg8rfHMhfgWT4
+8ajaEL/NqliFuPMSNFqoWlJG3fKUquNZrE7W6OMgDCiS1YUZ3ahjjBGAHw0MKGApeShpC2al9m0
mf1LJ4Ct16Ygko/H1Tv4VySgwZeVCu2ESLbKisDJW8gqQO5iDjZ6UZcbbeYcwjUcUVq56uUNL+z2
4/DnndrPxGr9A/0tpKP0I6xkzyg4FxFjUu2pCDEkRD/1uDyHm/9w70n1jN7nGQt13+t5Ca4APOJl
HixBPU2CbN7YGYdX2nJBq6OEXHKlBv/h3oT/V83sIrO+Yn2IcVhs8+jKMKMqI+6RPYK0IQ6Als/h
diO3hfWSghVQtJGJQf2J2NbtyqYVtLsUa8Gm7nX/jCKZUZbZgq2do3wuItM1wvMpRfBsRSA27lrC
xbnq8daS3j3+3kRbB52z+ItEgcwPRM6rGtwJpQ8VyevH9HLZpdfC/UKfTTYnB5Ge2KFcUSJkF6FX
hWH9GChqfb98eycRXrHnAtV/fi6Cn095k5UEcJ5iX9L+aCR1ItP1lvSHEjYIv5Z30zdWcAAy/JJZ
hjwwLM/QBT9JfzbH2I2XEUH8rkzijA7w9/LTT5nwvd7HraGU5ikWB8zIk6pUP+RCf8MSUWrjCoJP
mUvBNu9ZP0A01oJ7KjfeBfY+eUINy+TqK+PoxOydCDn74SkuWRSNyxlf/p0a12I0Tu1Y8yXAtk7J
niiHUaZjuoRh7FY8B1kC9vyvFyp1PBpekzcH13eZwD4N2DR7jkcRvvs5eXbOCgwiBpfsgXzqgPY1
I1e2zhQkQF4ht67xXP/GnADmBFyl9O5ZSt+N9a0FJ3t4EZnbzGkUUH+SdKyIPXTQQcVycN/nL7id
Hku8sx65+4u5mPw5yEJEyz0W7rJtqkkmJ7A0QZFHiLsSf2rXlGlCSwnursv8QGbPjQlUS4OQSuiq
VwtBnt5yUOMjrbN/sVtHc8BXK+YU1Lw9ahLAJSMnSvcosTJBvBX7jPyLSwbZNTi2qu1dyhSlRBBx
X4JaU3rdH8Nf3Bs2raNpN169Z3F5+kxPpZMPdchs37+2AXDzKhrNYV3yfWk6I2zMbkaPCqpozBHF
eA9vV2Yw7eFYZB/995Os/fBvZHAX3DtUUQCy7nn/Etuy3TJzqnMekme2Ef1Mr+KE1+CRXlrMSLsy
9RR4HedQ4MOfoAh61KDYl/VEEcU4ojNxa5WNyAfqQrGE5g7feW7BIT56JDCP2sw4TzvIWLC0foCF
w00ry9nB4TRl74MHNryF3xoQ/To3wQkaGdE8zchlEkVmVXVLVUc5OlTAhbTudu2bpOTo65LpWvvk
Tr7Fkx5/RDZ9sKOg2yG8ZhsOYJCOxFS56oRKylrXt3XhgJEj2yaKVnidvb9/YwFCFWhnLrfTNss7
M+h+LSuULv53cZvN0tQkIKPe1NbRT6PDNhpjjLAmeJacxqeUVsV7B1ZB3G12dLznhO+mr6SQQraw
+x+8rBCld6rOSNYFxdjqw9GKhkhcYpgcLMhwFNXtgrLdYZoe5G2b9Cw19lNIVK0HCu/Xq1GKaaou
j43fisCYREDRYht2Faee2RtY3F4IXN5iJkM6BA4eAQh9BSQwvqYzvpjFwqMomYEHqSklFj0nCOkT
xd1dxG7Y8LJgpWsita4l9flgyGELuyki1Pw7dkmekhGiGE66pqozlJIKxsOG6oWtK/qsraKXRl8I
sYWF8GAff5LTsQ3fkN1q6vySHpCpgs/0FvGPAVn1O+LbehIf6lZUAqhOr+K/cimz8/LtkaI4nprV
ODK/6zNhaokmS4yqQE+SM4bO6jYB7ITCrpb7lerMFhHcRyasCHapcgnsfOnu6bzOBcAbURgJg2Ez
k0V5rzarDYKKlcRg1zrYW46nU0gkLWzWbYL8G0J5o46cnsWN+d7qVM3v9b1hid+dJ7E9hOxdrDjZ
GuqGbtlzrIknXqV4FhTpKGz8s9654DolMGFnU5YDz4vy+mOj1HKbi3SA3aM72KZAeocdZWepY9NP
4q5DOqIcBOPhFsMGaGl76hERiNMXTcBCT6e2NJnTklSXTvrsa8QL5A18mzZpEMicPEqInLDmH5k1
fj121aGCMKG5mAUxFVDp0TrwxjS9hPpAo8me8XeiNJIUmgV1T7TQr1MB80JpqXeQGcq103I9IDw7
/Bf56llOKmlolE7TINPWD9CVzhNsr45NexNTJkGv9hsHROLP0T71VHPdET2Pw+0Bln3fbRiC8xFD
5qyozOJCqstZmxf5hT83XV8gEVK0TWawv6QLn9fJMXdSxuprY0zpnWghmYLTWpsZpRkbGIyquSNl
TLKsQy8R4sfxxerTNTU+kAGcLGCtfz92SAdN0onFx4sni6UNAfWR1nDKCVZAwk0vaxMhHHXgfk/s
RH9m0q9s1MNRs5W0l8Gd1hL9LbfYru1l417srCtkRCQEeSjyyVRFO6XT82U0i8pAejFyMDWOp8oP
/ZBQRnYBVyRN7nXQ9pQBLoMHcAmP8wwalyIHZNqs8QcQnpK/+dL8qu60KLIYYmE9CD7FxUVKY9Vb
PH+pf3EZW0wxy3qZOgWxbm4suiB3wMaBuuyF4T7vapz9f5SOmXDr/3kmvsLeshEPF4vBR71Q+UMs
rdnuB+YnQgJrb1+oR+m7og+Vh+oSbd+l+B4lE4mj09UA5IeUQjC9nOM+cNWvooo7eq9Ek21QNjxN
2vuYMu29wwq+UjRRW0EOnRLEoKHYQoZJyLnMG8iE0f7vTaSaFVtmM8UBxQcprlH4T8fK9cHUgwlr
OTw6+mnWEIPFyO5wiOSYpt2BU+F4MU+O2VmbzDWAOG6Ud2O8HCeP25RtFPpgvenGMC/Vc0QGKMbZ
xwFQ11qYWn1OEJ6/FaJE/Ihr1a70e8Ivlcs3GTrHarZI07yW71wkjuEkwRWYWtBrkeXJx9IcA0pW
NVzAcCpA3aBAwvXOP1kkq9Sc3jmF2gIUOO1CrUJINW0zXmxqxPgK9YbAdVqKz6ie70xxY57va5iy
YsAQ74POmzIL229xnRd7KpPAAwJSV1MUix+o1UD3qQahttLUL+cPgIECDPMjJJqSpvfZWZzFPfPo
AUrh5qGgc1ZQeBWIBQkEoxi+JjplpBQfMAkV16PFvaKB1gd/Lvx15rB1cdez7cHpNJ9iisAyQS2a
hSJLH6KJqcG7jzegMVZBU4EgaG3gJMaennyIBJjBhn19UB/OZZi5hHufVWrVn5o1e2smzLogVRTh
aaoqb7111/BB4eeqFLan6PsMgusdpZVp7PFhrP5m7pm4zvrteM0ttNecusjmsa5fGOYev+Q32OzE
mqdUSvMx/FEch4+dLnrTvUteWKuEP6ArdgNS1BPRKA+D10d11FbFmEzSxAoiuq77SGImC6/BHFQK
Xl0Ai9aWGLCN5X0Xau5uwtxSJiFlVjery5l591nZPJNJpHFZfxf6151kszi8nMjtpPrwHQdqM/D7
hQ9vSi5u8qhC4fhxcbK4lPL74Z+VXVm8Hea1ixPfQ7Zs165xIWkIpxy8GW4vwTEMShx9gQxcofwn
NsAUCQrsBIQqTG/+8kzsuBBtlbCIx+J9WA3st/V7b4CGJ3UH/h44LqCcl3+boTtP/efxX15XCiAH
7hUkyK47FAitL06AbaSh2l/Ja7QBKveX5+IMM8a1RfQ0Asnv1f1Xz6G9j1F16TJhxd6TKHyd5GK5
PjBKGWliT7TBC5oclVduR4+HAAoRF97YTRjKZWuX+c9HO/ZbWZLXqM7BbdAwe+ujKKetYFhStZ/0
yiS4BUqjxdbAhfISVIH+vaSQvFP3NsIPoamnQCfSnTYizle25h6bQn9AL1K7kClqC237wy3Zr5Dc
ISkob66wdQimPCg5PAU/mlsLelVqil9uPXAbF6h1hP4nZ5FMSta4gz7l6bNCBZVq48YHkp0O/fQn
AfO7nd3UPfInLDhgaOU4HFh/zHWBsZ5S5OMDS2DBPkv2/bwZYLMH/YmnISdhMR7r/pfOz4JF1IFh
WyoEbaRZF+2L84ehIOCENl+EMvxSQBwxJ8pmnL5DDUy0wY4mu0PEjEUKh6gdmH7MfqEwksz4943g
XPh88LCOgr4zX5412HUhJpIl2dAfoLCJgCNLW1GmOs6qk5cERV8PhYP2yi9G+k1Ptjq60OsFUhfn
wRjhu7Z9vnVUNvR3MVH/SIxDxK2kYGt1AmicfmCEYwPiES+iYcDrK8XT/IjWLuhwVgPXML6aqqpi
7R+/LmMoobThgKR7rbb0l2Jbgh619LjG+7afg0+DMJJTkSs44ta/km5RbiHPosJNvcd++PNtCDb4
8m1PAncUYdmzHCsO0OTmeu9xfe08Io+v6mVwXym2dJWPVubtmUvANi1npYsbdG/h4DbbS1ckoX9a
OKv4sod8TxkhbSCecWqk4eetinrv9fysUV+ZkRpua4E7QyLdxBcKogq2obXC/1ZpjuKfPV93mcGR
qjz5z07F/WGO0f6g78SKNJ3bcoKozcchrxZ33GrXi6lPwLePgdLfsNv+rMKudreymKTf1uJLB/ij
UupgztWcERNGcveaskLA1k5CadlOxH6iLH1Kas2pPgjgwxPJwKE6IKI5Y9L7OEtKHt1Iytop2aSc
7yby/W7b/w4UWCnVEcWWNQnbPUZ9wCuIrZ28NazueecZTe3246RBuzKwpIuxdVqS2G6EfFPyBtJc
u5c3G6bcBacMSR+rvL4Sqk8YbuyInJ+KpeSiCj2DsOjvxx9Uq/YUZh9DH+wrxfUtYgsXfPTUfPnn
r4tlUxJcE4xv2eUHVge3AQfNQmjcPfoFI+NGGqcXnz/NgpzOG3p2BfRy1YnT6Kkq32VRbdo7YibB
+PhSoSpLxuTnWkFhLp2lzyLayqe3qMoL3jPXLMw6rOpXnVNO8M2PxXAUWvx5Rv9WqgCIPtowbzOr
wjefFFHE01ajqzgz846RQaHPMxK2rMoXri/QOGaD3e6mPDYquvUqCoqxeFqbzadEEgJuO0F4oUT6
kst3Ba8hF3PubyzOiwvbQdJS5cILld5MNIbyKLtSIdhXUxPpQBTN9w/eB6cf2h5Xk8MQmXnagUEb
ndrnKhvDDwbodjjwQuPnMp5gZuEWw0c7Ry1C33mXCJ9OFn84DC2aN/4p0+aP5H2FdIu4FtJ4IbR3
5fsNI5TJF8A8NcZtjfCcBrVrJZdg9vCvS86fheDsr27B7c/EE4VhnxPBFj36bOjRmre9AeRfPyMM
dTeB1r1nkvCTXKzdJwkjVjfChb6ufex2wexQp5UkoXs2c2labBqZyCFg7eV0/iI+77KO2cmSx0mW
8S7n8hc9GXM0lgRHJ57PT+o9OwlThl3wosqpPs6jhUBPw+9W9uGM1fl30y28ROeFidPnqA0qCgxJ
jWU1C3iANzymfxWwIlcNu/Pshu3YVyj5nbuyngEkTOprKhEdB90fjxha9ishzXQfbvCArX8yTazw
SMj6Bm/opRn4etz0+PI607zdgXZJh7iC1w4oHzD7u+YaQ62oNtzrSvZtEjhBOfSc0EhOdkMrzOLH
5U24SzFRsekSKAdBXsXoS8mBMcoNB8pJ226oVeLs1faLM+A93LYPEKnpZTrsXNj5aZon0cAVLV/0
ml/jsrB2735UCOW1gqodYcF38E4fBTYWkmydjwJxVN0omVg5ATB/qCI7eC7eQHl5+yX9gqHwKPvk
kg+vho2jj0PVqA0LN4lyL03bMD5RO+EHdl1rX+n4CPDzX04+hBAU/MYwko5u+wvM/6DPzsXBeNYv
385/OpeuoFZkDBaUMfbEJxde5lA7TMuTrPm7lmdFUQLnwYxnP3309p93/vjBMLdI8fIFdia2JNqL
ugeuRO77nOQwal4wztjhF1vQBworJi7SYDsAacIQoNTjAU+NrGGhbqmpBAj9168zw+/3q4oKegTJ
/jmORzi7UnDdfj4X2lf9MS9rP2FxJ4QXn/e+VwKl8bTkul93FaMiOYF7H51bljG4KpghOd2b7dvM
DwGp7nxeGjf9OMr7UGJaJaK9ko9Riz/mgnicFIa5ZdN+2VtJD7quK5wq1WnwTkqlf5h0KmK7PDuP
Pd8OhlOxOGaOQq+FpyDyV6x55Arxnfr3CPvPKCUJzJTJIKQR9we6Htwg92OgEj/JnPakjADmPLbf
v0MDHi7KOoieO4u7tJN+7yqnstiEltu7yl9SGr+uR5TWtjfHEx/lCJAHvW0vz+Qqla+SwQzyXHlj
NqG7xOQwEdmQqUQCXzVh3XazrftChdIXR2lJiitjB5dy4qtWuBpRUu62l9a6uBC83kik31scpjA3
loZN5Jv7CjwzcOyoc+tj5HUVd1oFEdgv0ItAkoUvD4+CPK5dxROKKEUteQlOgQ16XNX9EDLaDhmM
uNlk4ImiSngSf0K7nuLZbUVntwkMNHifBxENJEursleKczMPSu1wTCeWKY0KK91myuMnMMOT00c7
gi6oTHE4FuZUBxx9ELLgHWdkfK146zymtPT1ZKyYWsY/xkLdAOEJDXdhLxJisLdpILsVmAIGLZ8A
hyjL409SLsLPsHG9lDovoMispMzcA3bfBAp7wq6IBK6GRteZFIZTcSQkqau8FoEj143+gS+WF8ZQ
KTJPQimasHxNTBOxd1yUkF9UeWlsziPVEGIELQw9UElFW7E/DgJaw12Qfv+Raq50oDpsFrEwdYpE
/R5KlmCS2wGJt18i5sHdU14m15BLzFOEBKhmbxvCbV4kxAhDqwHrkhlVDVDdStYIP9qcw9XH/AzP
RHRX52jJHtieFh4pO3zZTrPcO05ueXjnS7FshItvp9wPvraOda/zit06b2dslYDbJMr8MNxFeN/v
9S74inbRCfqTveg7BuWjiERR4ZZLEPU1y4p2oSYiuvreqc7DYDfJaE0DcYHUXFpiernb47EGBJwP
XUqfc0+uBmD83NyHF5mZGiDk4mlUJOngjorE4RJ3GfGnLJaufgBUr66t765L4nyPePXB+v/1Muur
Q09czt9m2eQPJ7813Um7rGqypE8F5fIaShtYc6Qd105QwmtoOprA2pCyLnn8vf5mM19b9FZi92Kj
XltAypDy+YE8sfekIRRqJqsz6X+6WdAdex8WliO+Qt6++myO/2ZIR2Q3SnAudKv2ysQYM/y9jnzm
H7xZvBBHuZHcLfeaq3hIGKxH0JcfaAaDFCu3Sy4Lm/QRnNLGPnx8W5WFJeTnhNeAxdHCtLM37qK4
Kwb5Gf/pI39AynDMtzOtj/1Y7drBVWZQQ+0A/zqByIciw5GswGKI8yCHxsLloiPVnM6X1kYJ/AS9
x3lJ+6nivFWbEOhRQQgT/CrRmsfk4XWd3Odok0f0SIcvdP1BmmgT6RMARrNm8LwJ8Lmu53JkUOjt
eGEhmyhmDGEJ+c6MyUdqIoH1TGppyzp/aSuHl3HJdS/cCdWrtqWrrLe+rcPbkV82/0fj7qLEqfB4
uHrjEQG9MAeIxlG4i/pRVMEjzSWOE+h5yVlIvz+gjRVn9sDeq2rPQriYhOrnQmcejS0nWZEYZ2mZ
7HTYhFMUhP63dWZyjVzdqCtCh92gbN+37d3e84eB1g7vFfX4zGGZj/tKJCmOD4LtmV0EcGwen/9U
F3RA1oHsm51GZ4lm0PrMNUNnTDEVvly3Q0XtmTZ5RKDb8KMSjuq1he3x2ba6sSquOspRTN5uezo6
U9ngMeCAc/hcay/bzxM4AaHk+trE5uW7v9s+vg2fXWq/UvnUGFb9NL/b5ETIN9yonDjwHwo79fsr
PV+DemCnrCyw8sO0KKBycPlQvcpSESa7dRiAM6MnmAp2Jze2UPTCZ+fW+/Ld5aY1J6T3o4cT7a0E
n0p2wkskD8y+EpLakA9Cahv2MeYzw8I08leRXwIjF+AlqSvZTaqTQ/jWWhfz9PyCSCLAQWHHCuY0
UU6AeqynQvZU3k5wk6GHDG5ZC1UJjT785JucNCVMcsI1lh7HEFKOUfrDFDOscHBEhXT0dGs309cQ
jg7tKLZgNfPn576QY9xcyQoGT8Z+q36FUKu/eHeSzMK0rteNtpi63mpccLuBc/wXYpGaC9dj9kQ5
mFu6ixktc0fDK7u9cwD6N8q/Q5cMsNI+g1ZqwuYysXxSaPNNYvL68M224uKWBmmKCzMVUFUCC+I3
7kYBLUUrdc+c9LADnbMKc4u3ad5ltXYb0OAFZfGuRyGK2yksNZfUEc+z0eCagN6AwSE2gX9tha9A
MJx74PZgXp3gmzn43ED/81RAGpWP2MnHOjMTqkA6knPEMgnTLtFB1e4jjw184BbLkORfihok0S5S
jRhMoXmOlwTXK0GfYTMo9qNFD/KqP8yq92zl1RBtqaacEbT72tZN0Xt8zzYGUP/9eNYwhHBgct/+
6GU+OPH/C0YJU5wfF+VMJeOXgGlymmBvMTYfMKhZd9FoyGL+wVqZvZtPdsG4ZTsk+/UFpbHh3jYJ
rgIhMvREz7WEJybYTKV5f1s6wYrKtnOOWRx2P1/RkR7CfGSjMsMYO2eNjGa9BmpXNRrPCm7VPngF
LAQN/KJSWRuLwQ7f83M/xt9jeEhzuoUZ449I09MDQpW+j9aKXuQYwYA2tGRAu9OzEYZrkL+YaBRw
nrpLHGES7+MYGgHSiL69qhVYLVyW+wZV7icH+WgESx58c4i+ub+2OXAFhEM+SdPRATRPV5daKRC6
xyenwDtMUU1uGkNV9/wmnJYFs0hbeCZ/CCUAYwJw7Fbw6E61j9b9aE4QhVEjs7xSTMXPLM4M1qAZ
J+TSIRo4M5bQItl4LCMFqux7Y7c//AonJNvg7KDNovb0tt05Ar2F255iDvP2kVvKYirHWInG0ION
E67Ir6fOyBxeHgd6b0vXdWwvoTK2dMinQof62E8bRbtrg4djAnYenjYa14YxGKXNHW4G2ATebKli
rNs96vwtE9MUXZqSDr8p0dbUsVfbmXjzPBlE1tOSPD2i0+dLHww3KsXSNu/ckNQUNtvD3S3MF7W9
8M5nR+S0m3ZOBnWwy1eMCe+5DKPbtYTnAhZanjjwmfyf2zoChPJm55zU2cb2sma7CVNPqWgqm4s4
IGy2PpfB1E+PPbBdoZjUhbpdT4MEQkceb7fqoePtP7uBVS8TzW/BQsETcNmDaQ+I3ucRhXdYdm9b
IgNt9YEltxt2QHqnaGeJYi5Du9RLaT64Cd2VMYavzYbeS1VzEvwiju8GFXfHoqMFafEp0EeP3eIo
jdt/0vQgud+7WzVAc4tQhFjDOSHCGIem96i5YzIL8hNYbzG9qffDst8qaQsd5kqLdiVJvNnc5av/
FCPoW67tTGnEEtRiuLL/ghTZKbPJkMNqADikMFJBicVO432E3h1WJxAOvK5nTJcVqcPoRYR3zqs/
X8x/+D+xAeViNdah0H85JxMFmrNrdsXwO2qX8LrnV8HPjoWZjovBQIH1iHHQi/ZkKQZeG2pT90yd
5n/X4Sx+qH2R20H9+onOHVPFRtQgdBTjar7wTcax5+NMw4SLbGltzqSUPxEJXD7bZ2mO674wIjEU
0YkKZulFuQO7i3SVfn0c6xmISBu6or9zdp1K84MapNLUxDEx8ruRDtYafC+ENnBLFX0+q4j8Jzjz
Z+nFvE13QnGSiLlx7T1kGifBF2HEegNW9SxJgCNdvqISmYoMxLTX8pBiWdBb6cs8KUPPaRvLqElc
l4bPOVwT/F1FlkNYCgLmoMTJMVXPfzWahFwghMbesCBWfgBzBDh+uahGBWwRgK1tyPBlGtrV9Wa3
BZKdvUC1i1C33r/I5kpRJ7khDF3qGi43zDdxoZD49nfZH+C3+/ZI3/Zn3en82AIjMRUJuawhySyj
IwyvkSUp4Ywtm76+vCWPn+fJk5tH8sB7SyO0tsnF9unU//OLO5+WkX+3yU4GlMATxRNY1gz4HG/s
vdwwU8wnkcePRu50KuNi4q5v2hBqHrBN4pzPSO+5/rHnNMxQS9/0DDqd/5qkDOyoNBvGRPdr4nFI
DZ5zfIxNSAqtfg2/AJrfpczgvZyzreuoODkqUgpRpPxxkKztVh8Ceow0lTyQmY20NTM9lB/MoIDJ
ST2mNJPuoiByU8ir5/uMyeJVaWpd4Ch1eJhJ/usNMVF62/361IVmHjD8QWPvH8E49zeoyEAI+8Ox
5ZCg0o46pXDLK7eJlUtGRUBGRtnheZ5W13vLF8oexfkk/LnR+dSiIJ68swPUKo4NJFt+bX/XRjkv
JKhTkRd9U8LK+3ss3GUBXEgtggmV6MHkhxE2TocTM1fZLy/LtI18goi1uGCA+tYp10L5v9jf6Pmq
loFvpEiLrfg5MiV7jqurWNxCBOqHnFg3LNnAQDeXAPjw7tqap5RXFDYX65/z05Yww5esvGw7oSg/
19o9QFe2DRWe7X7Z1WPTCfwG0YuwDVlsdKAZq2cneaQnTReE4J2eGVhClqM5/+YzZIWN+e0gx9R3
9FCPI+zpQ7MLZ1rM03331NggDjNGaQazdrM1W0fAGfpVhje4IrkAEAeizVqpF3fbpuON8x1Z88ui
NB3Fq6Yz54OMjlNn6c7IORovMomLvurqyyu5hxRDrvISV52q+0E6+XfBAc6TvSh1Q2Y4GX9jfmCN
Uc5oLAVymNG2zUHvr7AWLKDUXaw4MQd5u89BPbEfBVvx/b+ErVeIgMt7vQkcc0/JqbudNGkJ7zfd
VFc2P6waBbHkYwNWXuwIW5DYMAcRC0fKg2ZvnUVpzGaKSYJXRoDpjwgLuStoylIm9rKkbvKVK5uR
737Wwp1Efs41vSBtKrrAkkAR0ebmQVAjeCtXFN+QlmdYzcZbjM4pOGuQ7DrLcU6bmJX2jDM041uc
z4ZlOdNUqe05DRVGFFqVD2Fiwudb7TkkwocUqsD5ZaPQiLAPpjoTDT9HjkP7ERKOMKXUFFXpb8WQ
/gWbtgnFBH73F28ilZmv0XOzN709CiRo7nXnXrAgBDLDeGhwcquS/uBHs99xNRTuNGD6b9kJkRG2
XmnoZpNWdadKvnrAz61fpUq5qpAKCIBOMNC0JDp1B3LtI6A4fDCViuWmyKRm4BSr9bV8QrBZ/ABy
opadhncFW7wPHEaH+UoI8vMSaBM6vOYr1pLKvMdzitLfuUbJdN9ur1XUSZXqO+rIKvRJvx7guY5p
HDieBiZEmJ4q0WQLSkgDWnCG2pIAd6MTL0ElSzG8rQ52+6trzi23w4cf16BJ6DXlL8p+I+y/BdCl
yYBZl5dA1dJoQE3wims3sMxaBONZvkG+GwYX7s9YGm/9+lS7zcs8ivVCg8aI5t47DWFaBffa2N/y
2k6LDitB8uel59KPpCPP6Dnkz8ARsBhCgyvMLoPYP9MivwLIRc9Cg4iwNxBLfm/+vkvKE2+hFKP4
hGQsE9VlFT5jx6uDDtlsDFFllKk+3YOFB1K/v8k0E8YLDYjRIvODE2InIS3DMQa7RXSP4RzmQGox
IC6DsrDN+62dlTcQccZ1thD+rSRC7ZtQNce/IXEPnkypGiwBL69BABslrljErIWT/0RcTHfaRv8C
HXpG+JCjBQdd3Ef4gn/UcvjwjPo/fMnOa8az/cGg3tTMLXIUASZa1jNsetAjt8X2C1GxDhzcFQqP
55Dzh/rPhm2yPt/lVH3bRnS3o0Dhw8H81O4+IKxzJs5JKxzq280iZV+JITp5X73lTC8RXqGUbIYv
7nnLTsU0tYLGHEncvQrxo7FGrouoaJCPhIPhnMzOKlm2gL++k++ITZbyVBz9QFfRMeWx6H2AGY6M
1r5W1lnKoBbzvotJYOaIUdk5oWonQlZ511M0wRfbjj2p40UZGe7JyCkAJsVNl4llme6UrsYUWtJj
X2j7Q+rdWGL3/kAkbToKSMc9088wU5LtJvCy2jJJYW0X3Hl0Wypbygdpm2lRcsbRoMakdcTE9eCe
Pgs5RBNH0vhV62dEcKadtJCzZErA3MVVg6bTZ+c46tZmUy8gpRsCPi0jqajnAe87tJxDRt7W1hvK
Q/ayaxAoaie6GJc4LdRqc6yu4LeL59o7QA48DZPe7qBi0cfnO8eWFwV5cEBjBvavv3ddu0lCpDoX
IuWupNW7ZBN+Ej84p5zzbNqqVDx0IamRTHBJ4QTvkHc0dRwHoY8u0GHTRU3ynwkqUc4nRsHQQnMt
IleRqE1cr8SOvlEBhWP//gGlbfSkv9FQkyCmXI5innj59cV0fV4BfJBRKmL/sPiM+x9m1y0YeZp7
5rfnoiysMRJdWFyuXLaJok//5imXyXWlB3kiADDT/hVSf5/oyNSMK62BvUIGRWFKpFyPeg3yj6jH
J2jv0HSRnWvbD/rJW8QFAsToXmE5UDgaPIAsds0wgwmvoAcY/QnTy02RLNHfO0K+hGLLc2qMOInr
/m8tsOrMI5r/s+DwMu4QDZCZD7lCjKQNo1JHAsiKmg9nqDiMnB2WTV8Yzbib9/kq3eEHeEeo0UW1
1z1+0N0g3rfp85cBXRESbT+3nD/qk7+di/SQuR21+s3PRPxqm36BhG1dFjkNkWmJUGOkFUKOmFP7
BWVEDgolZFTL+ZAXQqeeXa6IATIjzeawVSDEpEhcW2N6EDPSeECJ1ovNpBFrC/ybHHzkxk514AIH
1R72FQFZ8NkUclz8ODOMYtIe46UtrcN0wB1wko1YF+StSAzWesLKKYoNKzk4yUKnUJEm0vbgrjb/
FF8YozZ+f5Z4G2P33yrtjCS49xrHkSeEBypYyVbMkMWixoiD1Z9kBtCiW196ORfy1Ee933QzZMvW
KV4Y0ZOdgjxxePP7cXdEq8+0DHlNuSzeBKgRVCPB8viHnOasqvlMYJmBqFBpTEm4vIfPYhAJzFU8
8eJpUn7hlEyTJ23OE0Pi9iU14ubGyDbKBEyU4XTxJ3xQnU/yNQpimoR+U0g40jjHGb+XGyX/Kwbs
gkYLCIF+PLudEU9/e5Bbn90AJFF8ewdy1V8vlFvFMQvOHdj5gnEc4QuKPT+flKNvOgKbAAQX799d
H7+iikDIsMq9VUZ9eQHi3AK+e+gGWcUIlGojQUSArgzJyYzJrqN2CBh1pKwujx1LoBs+EUMuAmd8
QBZPke53cPFJNOdUCeef2wpddRbd2nr147sOpqk2EHfqxILUooRCUCE+2jSnpmFxUgTNlcM3GIcA
3PUJ6Le3VSGeUAvxolqjnuTOS9JzB+6LrZmQIQVb5laMSR8mU3Pi8lwNwlFCV6SvzHB/0oBqimxh
fKGd3h6861dBm4kAr7W/KiiirhrpJeokch0A42eQJ7CGsR2jYyDdG6zJPCWNJ8pB1Dx17rR5foCY
5MVLBtu4FoznPrx1kU8KMOpNNppCHeruvneHVWyNBLII3hwEjwPSpUB3ConYCf3s7TN/R3R1FbKs
yMwmczXT6APG38V/SCHLgGD9t+JlotAAnrbHVpM69Mq+zhQMCegXAyOHKs1tUPIU1REgYSfeakb7
e6YSwL07c1s6rllwKI75E+Y59pNzRf2XUX4XJrxpQ55NuHBAFTpMwsAQBc8mOpryWArUuYCqn6x1
7iJWIZpCVRdVqrH/1LT9Z1/osoO7jzqGZ1kC3USPbTcX2Y785u7t14qcblaE0TxGAbcp+mq9yo8d
WdSoKCYGS/z1qoDBcdCld7Qzz7C/d54L7pYfrc6fCCCtI+VF/kAyE8DSVXWACbqFjck/j3bowomN
F4NlU84qm+Xq2CZ6bGV+oOR97fTw5o1jNDVlhg/tq7vtnPJ17YR32JLVwYc650qc1KTXN3xQeuUM
AxxWs993IQgU7cg7XAV62HivQjALCoY/QdistEsJq3hlnX2+kbNm888oyrDdbyfSSh3mN6QsgPkL
oXB7otPAgfeHgKTHwdkI+QZY+7Ew6FUiEZNMH8bAkyQM2apjXw7uRLjrqZUIkdEawe3gOl0pENDR
RiUHNH5nMdxbzaSwKsfPtTWOvApP7RSou/GICfFXGCvJqvePPKgQhVEUmvzwhKfEG4kt77i+uF3e
Vk/WsopLNW3WN2Wk5OQMG2rlYwY1L4rhfLdjhln6ojQZexf4ignzzzcXEqwjVoeJzsm0fsT/JD+f
tJkEDik7/XB3KuUjMuQMaQ/6SzLpXK7fMtlwk6ruv8oskzrl8fn3bbnEL6k0fbg7SzFu5C0Muo/T
78qkHdyQou+s/Q0C6B6KzAIHWhrx7QlS+sQ5f7GjRiYPCSI1zfhaoeSu0EPA0ViqgzVMLpmWZ7FY
6KOLSs4WpzGnNGTOVxF4YNg62qhunCrY6ujuZt0iD+hUvXlO+PiIBFC0oerc0rH+VZ+F7y6TbGxw
8kuvgSQ5WG/tGEq+wCm812jfew2ta1DakVs+I237Q8HDeMdBFjR/gbXd9ZuSJbw6Z3fED2tg5B1U
g/byZOz4NHmBBI4uE4TDND+7GYHAAFOFDZkbGAZt41C6bKT8FsP/kbS0ENRMK7JOlf9nDkQVCSYZ
bzv/0IiKJAEILCYfElXcTpryyqDAxG0OTL6rIFWF594uPtJ7YeyV/nG6eVttnTm1FhOkfWqA/nUN
749AROJz4+Wwvcn1q+VgpMdkZOKnMZ+hnpEZg0F2daUs+P2tO9kO9/qGZBWXBh0C3kJZA7kThKVn
apdoZgD5iSCxxRYqoZ8I1WFUFHCAUj4GPmpwdYjb0FBBCjBZLGz0gMzP5jy6HdrzgRfP93sTBN8N
FzfwI1LETwtGPKoZZ2GoMULVrH+vQQ4kArdkcWX6kMMYhgHuz7//hhllsqdtD7DweBIH7weHenx6
Elf5oDaXS08fYhRKqIdmEpxXujKBgfAWEBwWW86acv6WuxxytOU1HYXeGiTDqqy7tuaGX423Shsy
/w1HBF5bG+ub/Oq/2yGqaf0PBAmns3nNI5CetZhqZf4rWSKtlyomXICWdrTfMnlZDqRhY+5XFHRn
Q6wwOx5FXzEh8HbE/wgLyWoyJ5vhvDF7VCCYFv0CUrqhIyfKsDg8Kxms1seCJuXMCCqgrn3PrfYC
8gRXIdzncSjOHwLY/vHJIz5CsyJaozBLg/6aundela1eGLdJ6jP9ung0C0svjRktKRfzQIjKPEgL
wr+an57I2wTHo7iQ5M/810/4W164AQUrnZgq3uB5tFMkAU/9q8b8DhGpuKLfiKQNuVUvIEnMVKFx
M8rTPfVGNPCLUxrC4hyjnitiGx6fcn0V1h0lYJLfQvISysEw1DL+nGX8MpYoWJM7u2ZoEfZwTR+7
CIT9R32rbKsDSEbRmRyPQJUZjdGctrJVd8AIuBP9vUTnfAQGe7hiqspHeWvieTPAFDaeoip3zA2L
PoNCrX50U9xU3uHq3CXk+Maj9YsyinWqxzB4rF0dtLcmoRVJEl4RBClQ5WXh9zlQIJ3ZofoYzEcZ
hy52UOBmE3QOZXzF6xNGScY5jRSqedpnX6ekeIyXmjqShgY0qudM5dztkbDRV9NaLCmHbC7FCKll
n9u/FiOL29jjDGZUvKixpAhtqDTIvFJ3yZ34gSP+pfE5/bf1YmB/Fta/+txk8J9kJ/Jv7QbQFpLS
O6k2QKGURz3PTL1D7O8No+HKD3j4qeUS9I5c/rQsTsS3jldvqP2S0XFI1ta6mYNVA0v9D0JHF/Cj
YeiDzgGUYQ8HGUsew8O3cNwnB+fPpWG3RyFOQUkuyLiy/SLS92AJUMQGdM3FaLBplSg5vcwzVwkL
VxddvLsZnoR80YvBjjL99y9Y7PS44ZKc3Jat1yMToNJPta8AUs9vW8qGRpimsiiOcH46npqBERaI
AtzbSuHECWrmTUIqXd2daM8Stuu3/xcckVFLRYSBw9gcbNLQ5hgsaSjqEiP4Y+IE/MilERF6CuPH
xMuKXtJVsuXWCv95Az1onIOjPLvmWwXmP8OdSD1dP/d5IiO3H3VOzn4ZKWHY3dJyOTl/oMG/k4ve
b553dysOgDIfa690fJ4SFxj+Cjhc3cnyjqkv5QN2D94GqUMnDx48vKFrOTKtX2ZfgnaoeOItmuJi
DTo5J6+6PdS1wXOLAvihlVgCe2cgF3hySyRmf0jaL7sYfuIAeHYeFNrgRKO9dkrN/zpgEIhwdkfp
qUmsQGVE98caSGmnYrRiyQHzjWcEHdQczb2jmsa8knKi+L/35VRxUkM5DgcnK4k4NOJ5GdVMbyu/
55JG3DB6/YbYIjTbnBKuOLMDF1EY/ZEXL0/lKtEtTJcCmYKSsBnmQ+Zsn3Aug7Vi8LeTvug1v4Vn
edZaDuIEBw73FagLQvj8SSYwVpzX6NzP3LExK/xxX/9C67WiQsDHR95zH4ojS/nBiY7Thc9cuxX5
kPRCm3u2Mo98fT4Is/aMuZ+0iB7ii5gLMZWLPVyAfGbpd8MKw728rmF/bBLuwychjup/qkZZ0IF/
zEWPZRatjKg0C2cMGlpblsuDOUhmyRJfF+2lLtvUVH2A5mVXyhmOTslNOUcbHZhQtfA8HkvF6Pq9
nBOHQRinGYuuJ+Y+XY73yx0rFgK5pQb6uTkWLLSJeCiMmKaED5gxLwOizK3C6tzmWnLCh4Q5gJcQ
F8nBxpi0FqAM0jHesg0rfcJnjk6GeOibk5cz/+wZhKBbDugh2zCUjBZpPngCYer/jhpVBCeFDT9t
zFOoo6aUvudbIt3SqKtdbiTE85z7+E19Mxs5+IQx8jVZfQUzmMOuKfWS29k3led+pKgZpgCNjpXC
yeEbOeg5PviNUDWUweQamv9+f5yxnBxp7Qe1b42U7qDttRYFWmLhy7aqXP2/IyVduJQk+x9pGqFZ
nDT/hxA73L590npQAXBY0SvDuMg2OYSUQxZAiafNWJYuKLDaZwTtMHrWtbkzragrx2QYYeyUNNEw
dPssL/Yxtiz/ofwgWQhIA45RwFlJBjnBSXmaOqc3sP88cKgLCXoBdDsedsdnH6rokcqMUaN6fJ9c
KtYWHONmOahgZhCT9zR8bM+lk7iC6rlr2dLXtWDrbv80wpC9jegVMBcUA9hJYb//QVRBJKgeNDjb
fy+ADNVhu8Arx2FBfDjeDl07C0CbcJoxQgLy/n0ESxe+ENax0WS3C6vt9WMNUeK7x8Cg3BZg9rgb
5inp+et0I1ExS3e5CdL24JFKf/QULk8oiMrdkyGWI0HP4K+DbYOvTz3peYsdMc6X6IBiCJQX3K0j
uzKIcNbYjcjJLFgSY88ud3pf8iGjRh/R24ck8zN0oIaFaUqVVFyhJC+v6fYKmdXjRUO42Xs6Vo4R
kVhaiFjOY4Uq7/NCiHOgqhLr894BmttIZ/DAZl2DOluFtXi2GdY510j1Bm/l36QEDnCUnaYHUi9F
vud2kc/NKdakpzeugCZMe1mYek44FB7NgmLZOc5aKc4+VY76yi1nsOefbxTS3z4FgV/0nUL1lD+3
51s2wP9KEUJsCrapfxSftASdLh5TBANUz6yMyABre0Bklx1OlQaNvU86S6onMeHyY/cMRZle8l80
8jvls/TsSJQotbMLvJB5R/YpaOYjHNGAGc1zTHSmbLujLccNM/UaQqsIKOgp3KL2TSztM3HECnzj
BleV6aLqBcJHy9occymG0NcvUSY/KI6ik+CYVVHrWN9vAt3JsEQyRxbRINMbqbHuheff+hSNa0KO
dj0xogQ3Cyc+amYg/yZ13jICfquFIDbp95AfXTaYoulVOenDkswQzZceroe/ICVynMZ4XCNRiIxQ
tI6yI9AsQJbdaMPS9wk4FaMEpiuf5vliGkXoObXI6bEpdTqF2REWkTUPlnyS9wnzGpj1ZrXjbgw6
TeIFslbWkMHCp+ohaHaB8cQaxMgZBsDzBxIpegvbwS3GZVzO6LA1n0GNXm3mLYyRUKWnHADKLpd0
eDOxEkxxxFKWTiahwvlfVY/Xel2r5NuzibJhsJCUH4/buFA9I3YAO43SvyCqd4te/mhW7aHi7Tha
GWiI+cnw46Logb63eLedkDYzS+azpDzNZu15l/FndkVNbVYVXHikuPaS7wCGwvVgfEVC4ih0RMIq
ABThFqwuMelh3z+1YCJPlZM8KcvNioVAh5zSNLdjipeEF9EDJXiZG6u3xePYc9GE72hSul9cvNVf
Jmscf74WCXFtUlaHfAdEpNPkwDLmqwpONsUPQ3zSQuf7zsxdQY+EqBqZWx0nXVkgnIAX0/nI8xVv
yUCYNW83yElXrSfVLn0HS6whXGb5aqc3+Nk8Ou0nGOHQZD9ML1GGt/uQfzKrv/VhYPX+il3sInqw
1ny7SHohzPaMp/kPkqmEOF0ioCePARCcXDGNzARNULWWeO6uHw2+K/suKHJKl9/8tlmUOl09eHT0
DLD1MrLdAR9aHK9IjW6vmqphqJsP5kYM7IDJHyyoS/G547cWFmqk6txBvBPc5gatjxbiIW75QPTa
7j+VmTs5K/9TSbCgyY2sFJrabExqKfUbN+TLWZJQ9fGHWipHNqmSb+CIgpVKb3vO8ND2Bwj+MRc/
YoogyX0hSs4t/IrEQUl/Z+uZKjZ0Eny3lfQNYQ/7cm/rfROuCrJrkwTuvpj7nrnSKZxZ7cido+Ra
YacnpuTasA7ctcZJ5tDGCkpz+o8wvKxqvZAgrNiSWd5OlxoPLotlkv7Cg+zXFMnPIeeO1Q98AdQA
yiGr+9vCbGia62M2sEH7ifmOMCQtynDXuLyHp6rSBnTnyyA2BgivXHOFyAeXkpRj05NlvtiQ/kIe
hZF0jhsacxTKB4APjDAeapbaSl6gyURzHlDhilm5tHMtR0CjuM5UiG6FL02fyuEVbfGVCyb68v9o
owOnjxmIQpuE83rj9APpFN7XO1SSIdfusVHUUVKcnGLG1+tdu3QH9MI3BXZjNLP8XilZ7EUpmgPu
wg/pzV+uFZaIWF+98ndtNfp8pxN2h9EmNYscAe9VSTHmTHuXaAuhgf5yelEya+xCoATYQoP8SVkD
3KDMEIPz4h2JP991W8za6zNitmE12ml1UC/FTcNvXWJ0wBek+yaANES8ZVS1YEzrMly5UtsBoe4a
JjkJGMrumef9meLOca2H93AW7Wb/u+WvXvcrNb1e/Mj5oCIOESnb6yDXGK3ZpOdfS1sEr/ftD2tr
r3RBNWSo//v8gbyE4vVKXbjWmmWLeN/MObAAwy7IQRsNstpXcbwfMPDECHBR1lewVjN2dwG8gZHT
xsgNNproAPNV0Zm/p1Pc88xCgxnai+JSu0NhnK8EJxgY3c2Dx7UvjeTHYPKUgYXQ6n7IZBqJgZC6
Lm19Ipf7gty4rGt1zwWVdX2LwmoiMDsOKRoGY5oTpBOQDaLAqMNSq7HdM2cv5UuUiQAkGvWJQzUy
1/CTgEr6FL3outPFMUVWaMy9aS51ar6rMyL0JzqqZQjrecFoUrCVRhaq2A5dxYhj9Phf+KKKVoKa
dIWwc0bb5XpMEMXlDCJ0MYEFGm+XGvv1kXjXcRYTo7nKNZ4sYRpCaHRPoXxbp430Kvjx61LXB4xh
NAgTFQOB6JfQlS0n99mae+mFv4Tmbsu/ZTXX9EKrjBS0HBSKh1OXa+FkAzux2G0tPXPvwSXuhTfS
gM+ZrECp79h5N1YHQ1PzPVS4uUpc6s44pxsr8DiVm96l0783QQqwRm5ZbYcjiY3X2OL8/Ed6SzK+
cpZdbyI0YLmQx7iOB4KDSJLw4U74eqvp1x8o+kf3G60iln7Y5sOhoPmEb5ExTXLg9ZEXAhHct1J9
KV953RG3R/k9tkNIk/6ZGY1FnryN4Bv6hqMbKsaCywLHKJZa9blY1+dFcrzXoMffaleiir+9GAZ3
sAfetYvR10+Fewkv5k2ltMggcQ2SuylEyffxDJEMojwJxslWLo34MMv1H86j3SJeFZuZPq21tuC3
69QK0nAWHUBDPfhjcZjxMTPJbzrDFoJAB82WuV9JYVG+ATZO+rMa0RScp/Mjuq9cHtdFqwGgXjTe
XP84qEiyIW/qU3duX/OmhasiALqDPRPIPnED+SVOQpByJibka3mA7CKl1x3Jc3TIeUYNeMnApsy9
VIDXTWpCFFCk3Xx+PGfNoDQ+moxPktcajm0BWYtUdmJrKrDIjRtAQatzHgzBTWK1Il5fyrr7yi2O
EdaDyGPHJ2yyGehCS3kYHnvVIDCAdqoIMsiOPMxbZ3eI8is9pBMbFWKY0PX7NfRwgroAWJBNF9Wk
5j2Yc/57dAZAlmALqGtP8XAepJzE6C7yRqEBNolPHM2PYXuLjvcccvagTgRnCoXyjnxvswpSho8Z
bQYfXzt9KywQ02UJUtcQ38I48fZX6kLbdsmyq1LxRH9xrkijMFptN7jqtWTGNbYzYQzcDtosTSSi
43LoHl4qPsIkQ8B82IeVx/7PL95xNl7jY0H1SF9unNv2DwQDFMMqhExBi0K0TuBxJ+ZsfyKjkG91
1Ma6Hk42D7vwbB8rLO4Z3hLLzUq2VB2IlLbvExIQMbt8DkqbWLjo/xtUOlt0Lj/0Gm9Jz4SooOr6
MnpQBMUg/n8Us0fsDwNjhWtn9oi0MS5QPkhvBObCm0xWUpTCgK92PpPFGANyy2Y7Yl9AIRPEIp+r
UCxX9Gk6qLO6G/UzOP+vCdGZ4rDlUYIZuBWM/z0T0l5dQwOlRSM7FXb1HQMvrgRbp3wUSgyOkvWi
cjtYXowMIOgA9nlrBDE/oLHObpjFUqyg0K6lBaVmguN2/udTVJg94SiI11MMdevmSjMR+ov2IKl3
P5wZ7x8cScbessgZjewfrjr4HSjL0R9ZdAZpbHvEkgbMA5RVOG+yfFVQGfepGBWSu7kDwwTP3Phh
YY+6RUpSnm6PjFboeov8s6kOi75Z5/le08iTcSxOCXyPMEUG06SUzsbZJ93hy4PWLN46hAmdiFKC
up3KUDDZcn+uoMfTmwO9zaBxERo4zLnebMZhIh+pcKBqY54Eqp2Da36pMueOsa8Nh26CZK+P6a3n
HIuHVr4/f5FlfavCP8oSUGZqy2Q5MNwxc1w8u2BKnrOISDNFxUmPxqeGLBYJ5E3o57b1jPWb6xOr
Zg1Fw3LMQy/dfOGG38TVjHiqiasF0DVKc2368YVoWcySO4gDAijD7o2scON8hg2iTTnJrfrV8Jkz
tRzz1LSi4hHZduUtlrN3ySk4fyPfi0paoToX/O5cX9h6kOq2dVIC7jb0cTKZKHnripyrZGLTdQMD
nGcx1J78VLcDPCrBV1yBJnWd4J4nH4L+3UsLLOJQtfZVmlfhmMtx0SC0SgZJ7X/AAxhiA7EanQYj
SGqjw9XD20IFQasBxHvZ/6CkzNuLQboJo18CWgYN6RjYMVITcm6EVFavM4HlCt4nlwFBulHlqHIB
uK5E7ZK2EteZx6PBAMfDVkRc/KB3LhZe4S2x+rZhwdRk75WlDFEwxozX8htcnOe2oJk2mPDpFA4P
nvGkeBWR3QdVll21nAE6pczZj0TQjE1AFTZVeHDQUEDGsLEAXQQV5Vt450JxPiV5AwXv/450qOc5
6rzEiWGZkwCUz9pWpVkjX4F/DXk+AE47Y97jzcnJqFW3cmU1H+1K09h5z9B6GMD8fmcTrsKoLCVP
M85g6h/JaBTX+oNuUJAJPW/tEoJNGqUUhJ2KQ7Rei2cfeJdqUAi1v1TLtYLF/mcsCMS0eh6VY3ll
rGwvzIjffVwSYCDgtTCP/gGGCMhkLBRaa/1SqR8RN6BbREFE98CBkaFA4weHKMUR3gwrnlUVtDQn
wWy8NAt6rgSocMV7SXCdzdeFKYRm548OtzbcLUqyVZ3T5lEbKW8cDvhHxWVnH8MihkqdYrXDydpX
busW3JXUs/59vwKr4o8TUoNvVOWrOP90VODFmBUNkMtkflN3XC8C4qWMgcjgE2ggwYU3+4IXKGJF
DrB8fcs6KowV5kwEnc4UFuoxeJ7AzsHwXBWyyH6+V+v4WWPF7XfcHq1kCxD5mCufW71pXqszImWa
hShSj99tjC13/IQ3sxNhoFsKO0IYfC1W92W27cxa7sReYzLQrU6o4aiVRxCB82egd419/niRSBC6
PR/1amfYXcQEtb6fM67grWGhXF9CMZvTXBdgfIQsQnuemt8rm7mcim0QV3XoreIJjWHwU70IXSUb
dseuh6pqvS079PyLXTpdPaq+bikDE+jbOQwmUwMEynsoWumxffAFaiHpek6ixPwB7budVQ1+O5Ag
muGtS1EFEqPTgjx9fauab5YrcrKEym6UwYIOgI+ymOYQvxnqMuxtQ+ujY/4LcF7xJEElcYENmhyt
KWi7u2e6IHmQ72uqEc9GNwLC8561+G2/yOrS/kvwUPEtIPUOxPOZQRpfnKS2F7VuhlfynBWd7I0e
lqRvUZG329Ao/f/h6TqTzITCLZZvmOh4AUuqv24uu1zbGHXy7DmqrBc81YGl0wJ3S67YS7mH3Xri
zRmDMIJ8jPDZCoCtd1RQJQvALsxfM6IVjUuFdokysauwNWgyGkIpcpM5RlVGHzYTQbuaQlqeKC75
Oh+U3/Jg8VK/j4uf+7J5p3Qos9Jx4RLkLniTgHsYM8Seh59nbW4JMxvQqJKcXV0qWWCTrKUAYLIp
afWSzxq6zXyeSvg9o5pWGGoSB/ZMIO4AmuY55+PbAqIL+vp634sxc+rbeZCNLFWKYXf6iLQj0iQP
tcK9ocoFSlCqe+LesrmDbyyasv1IH2Y7MH/ns6rFhch0OgnXCGiX+yIRQawYc2LmRoBCWgRTxRlB
fS5AnzC8Z1rncenoo57ugBcvRJo+O+fqsMkgN9aznpeJUi7tqFFIENIBOhb5w/hhyNEvb07Zxo5B
Wc+zy21m3MyBWumRj6ewmhEoC5v830FHc3UmBNXUnFddBtONb0T6lor3+lG+om3m6fwo0QB2rCOW
tkVaC9KlPX2W/BSSGJYf6ryjTgSRxjanf7UP/g2EUAQN601yya50vMjkouqRWijUs4srI9alslY9
u7YsJHStM1brsjExS6jXI+KNRSw8C++z4DiFHALtY83zFoVh+csRyC80cbVEEFS8qtsmIstRpngf
pt88YykWgjpDViZYeOKLUA3BmwRVfct2C+yV8KXORZAZ/UagiyZvih/FaemhJCaI9aLxVt79qoNg
0DsXDUvsg9GcLiswsnVuSe2m+uLquS6qsBbfoNBPTAc8/IFLxGUJxIB9CS3wMM+CPp5ElMILz3dQ
jr3nQVhCvfacJv0CSyv2cUVWoTHIRuACvbihhnz3I0ih15GKBXAPDhecntRWgtjPD1HfV2AiQuc+
2S/dNF/3dKSqGt4avHpw1RMXOidnpDD0wEzU/FCqzalYXy/qKQJPfF54hKSV+USOubAvKqEcQrwh
xH6r4LV/uP7wjxZtPwHfcsOvYK0nJaCnHkpWv2rtCb6tl4bHDY6zo09r8iOfAiuh4zA53fTPcMPx
r7mc/PhIOn64yNSGZxK9Tghqy+JuvZM3VrBz0JVZ/lzsPI9JoMENc8AqLwOUEO4dH4BdsOp+Pe7h
PmFB/JUYmpIopIHaZlZdL1vPMcKX8fW+i30FRkSorXy0YCdmhHegpC9VPvptyF4LE4hGoCJJ28hL
aIzjh8YfY4i7xcLmY1FZrh8j8jvnoEDiyklSf+7WY4VvUgZnBETjLZxy6evIlrojkKyzAcv5z2/u
yZTyQ1thVJxt9Y+bdTChSPSqUydCBtf668YDV1dMxYtAqLB83nDS/om9VaQ1U+qzlt03ZiE5mSuk
qYzc1yGKTR6RM47V5TV1lcatoBd3WYRfn32K9MYURxMZwkjhoshv6zGKG/b388FWoghz5akcBSeh
cnTVi6TQ98ItNlpFaoPhdFA8sSI784fSF9yGUeNb3OPhEMXKyqnwU9E7gzymkT0BqmLP2KjU+SpM
1wEAkjjMDPd/cYhvz7HFO+Knv4ibPlyTPyn/9bq9gFvAG/w0P4+9aUCVMZlJqw+ATPoBka1t9zBI
216hvLxKx0WUZnc59PAZE9HkHn4BZ4vnR3qyj7kU/AX5cICYFXFXdKP92Vystj8Yl2Yeg06ayQyO
ZXXYImpm8old0ISKnn+TF+glYAQLaL63wG2o+fpN5JPU09zda3sjtwiHOGqDWDM+6ga0VLh7MdIo
2FF3Q3ippGxR5Ajoe/0f9tJ5IwE/QgLtqD6EqnWGL7rin7rn5BndHgjSntwoGpm0s6XAx/8OECh0
iCbNy7f5YNuvEo4nBtVvPjuLVbTrERIvmTsyxmleFLi6ZtU/Mu62/+dYzArL2J742gBLyr9wqAM/
w/+y4So1lp2k8ASgLDvz83UtbAs23hv4hnBgFEgUrIkugPpHOA9AaaxJ7RaD0rbvNlPKFBF1p2UO
dS61la7RLo7bePhjZBkaPj4Vw99UwSyvP8USEEkcmsUUTg4tJvtiwFkAW/ZNfTku0WMHBeloS2vR
QBs1r21xnE8jBQV5q92daSf9uy2IvvaxcczvJQli0YRpSnTgILmb+WUCTZkRhtxaB7ykEsXiQXag
0a19bvfKmTPlbTQ3+opAIBLE/plFdwYx5y/dLVxtn0opveBU6LFKsP/d9AbBjvfBf9Xwdioenes1
BHw236CR7tDsBQZWVwb3FoK7DZ2lk/QFIsteEGkgb1sO+YP80pYW4jsCl2fZpWL9zAr7bKvFdS14
guBAgViaPO+qu2uvVB8XHLbCL3aPcBVC6X5uD7x9Bix2xH1c3+X+T5Je0nnai70T32uE4PgrVYVD
IcyN0bjenb7bpi3kYoAVl4oFMNfeA/7J36R6YeUtdCbSheaFbcfyv9KfT5S3Iu42wsHVvaybloMV
dRXAGfls3WSULMpnyj6ABBGVXlTOddtqYNa1kPJh39uYTcUx+j0knYmXpuLDyTCExXDyhn+N/J9T
F5SW4zG1cYjuoOrRYJ3NuZvWbytnau7ih+rN53Qgb28BRjL3v2oxgrA07TXLYg3pGNp+uEh2PQco
P7lY87V4/3v10fQbx8YTBr1xqjghVqCEg6XXJaRUVIR+x6Rf0sjPHexczGdmjtf9qOyEpzfEo+Cq
QA5M5uLiI8diZV5Bc/XeFqphcLzubMUxAO/T1CAxdEaBNZyO/Tow/V1xXw8dL0N0IV4OJZuUxZlU
GjTEM5ONXF42F8IarkbNk+ftr+6aoInTPKXfpeLlHGs8Bp508cXzvGXpxdIcQbcPwJQs3oj4cleI
wkgdbr5aeLZSn40Xwr5X1nNFUB3TyxSnWrLfMmbrV2Y8KOv9iLNFjW9KEQUTFwVt/O//dMVMT9jZ
LrmAn+94V69SyWQOeMic/WHP9xvQxWUQfF2ZVq0sXDpdGRprxWURd+zgZlVGtIBvIB5mUONpdHPY
1m3aEfAWbA88TNu5z6iZJHiAFq705fG9mYcV+5BHjhuxldB9EMKsg6oVQ9VUeLrui6iRaUDubtd8
ld1UxYjDzZ/vmP70oLA5ED1gVHgGFhdm7so2VKEY+BwcsGy9V2XOBKrI13/p2ZAIY+o1VI38wzrA
f7PkXISPULO/o3XKmOvjBEe8OEMBy2RhE430fglvaWAsZf7rALu5MUboSCeSTTSTGcsmfptIwQcM
xY/06Tyo1pBWqKyVJTdalQtElHe1IIO1XtuVGt5SGwD+lJSs8y8xuTYNiN6gYVoHuae+OSRpC7vL
t5vqk1DndRwRYps5oI37bso+0OJYbIsGlP4MxvoIYYxAeMg0jaN1qRNCsQr1kif5bmhVUgX2tpY5
xGYDWVjeDfk+9twh4w/EcNeJvtYocw6SmJXQVIlgEKUVlWxXh7SdnpeK8fJf+PmeH21VrKB3dcvm
gniCzCZTxLivOpImOaBkfOmoPzX1lNgwvjkqL17Qzw39aiWRYfFDETfJ7qhPtbgGz7Vm+t/ap4f/
HrNdvF4uHPnrg3slPvqjGkpxTZZV2VvIBAGto53kZJJ7pPBVCQtyKvLBU931TUEApZBm7JdzwRuc
ozrgXmJpdIbobtCxdpvo5pgq6tmYvr3C3si4UQ46ZMVlmjj19fJv8svAEUfvHvSAtsX6JWpDWk0v
AwpmoWXra389PJgNt5wdbRnziE7L/t/VgVVCiyzLbnkakjzW/24R0S0/dna96d2bCgyDHaKLZY/R
LLqgBJcoJs9DBYucLNik7mqQFpdDPHBz+wJdd+KT0HusbrVTrsXnbpLc7akTvWF5YAcoHO7pt5zh
COJoRNWrfs3tS8YJezAFVVTEn3suoDmbWsxSWKKs3fBLwj8mipqJVTTubtSJ4knHQ5xYdecNxYr1
R6GQd3I5lBRDCCwDRljmZSzdpckOHCo2clKWfkzIokOQPC9v40bG7GGARka5F0sChAsuf3X8nkTg
F+3be+3wVzXGmnpDfa++Zen+asrRvpyvKzSedL5yz3vcQ1GI/wi47iwkkTZg1UKpS7SaD5jmNxfQ
gHqvwUCeQ2Xy4sGcWoqvOpp45mO3hbDnudgRXEkb217EjPOA7OHqsVUCLlOcAev6DeaL2OFxQozt
zJ80ESdr1ZAA5U+k1LB77MrhEAeAiX/DH2ue03sRgc1WzeVQ1bLo5uBFRO8E5XgFMdNjwF2+4SyQ
CXJCcO87jFpxAZWe4eHjSlldDlfwIW8ycoAiCE5Bb1aIaIhS6a2kqbrSHWtztWLV7qGWIIgepwIY
afx1aCM7QCs2f70XxyrDnYYo57PX/uD9sfWo1qrfUYrzRffQLK+wGSwdPYNmnddvYa1vGoiee0bQ
vMXugtIPRpTZ1POHa4xLRyF2n17CndHdpELAF37uvo1db7Vke9XHrQT011W8lL0o0IY9CqodcZdw
TRbjKHg9NWRGOLhWBrrEzxhemP6Q8s66D0e2ALFS9m8fI4BUwMp0dProne3GVRu7zkeZRXOJ0vj6
6h2Rvi2jfzScDucJ1/uNrXRnmmJLKFhxHvNWjZhl5RG8BPSfGZ/tCK5m7kdqhkfkkeUP++mxM3F5
CZFAlvFr1Rk1IkBX+KSJvajx2MQ5EajtsFFfVKU/zzZV43qgeLmhDtZzG8Py3Zx8icb0wlACnTvi
WrUXbvMNs9TEJu2EcL7yP2GfM3PrUlSyP1jZ2oxOjOfy6Pf1cxMad/bTSuJvX9tw8g3H0IPiQVnW
3do9Nz/QLuFwWT5Z+yDQH8Qc+zoLW/3JfMBffcVnw3FfghM7NGqGWzWPrLEl048Tl96OFdiwFlqX
rnB8qq37GkhYo12SYH3SO2MxCH00ej1EpaD2lWda9jhKvHEuIfe3ZgPt+c6ZIJ7PRhzJF4Xvaxn3
NI0IUoZVGFAjVHrFWleYnBwikviMg62/zWOJX9DzOnvvJr615I6b96t6zp1Pxd19FICDRbUdGmhU
dxwAJoAW3AtGubSz5Wt/ICHuX5BNMMBqIHhqETAi2NhsirBUvuxB9g9S8aqrwggYvElbitMOb0La
v00gtFMRqbLgMRhiBjqAD7ac/VtDQMqapcRTYA9Zg3OnbsDGffPnxiA+UMobHG1OKg5iNyBniSMc
fVfdrNNTRBqcbFVPcH9rtUujKYhzcIUAZxCpfb47WC4noQA4hOq8+Z0DNbtgTvcGfV6Unacoz4pq
/i7BK9pnvrENFYoIpaivHaMIjOoenY7Jbh7wEpliS5Pt6HJaAS1SvujHonvNyVIPDVp+MImD4k1f
5SDUUFkA7TdFQcO6DSPGOkydrXBxZsxy4gWhqGk0yxObDotElFLeKJlv4pYRSzGL+ff4xaES2+51
rz7PKEZt71e4ci0iONWWWe8a6fRkDvw0IZ8oH7R6Oc76nEuLqheMvmYIhPAOL6LvA4wGDZkfpMcW
Mu1VH7ZitGBfadaC0HiCp5sXZY0+jseYfdK7jpBupEITzcuEEqCv8Vcbab7TMdjx7YA37+6aUkX5
8GVyqOiLuG+xgYMkQx28FEIEOMro2svFzpLq4Rpz8y/y5b0HhrfRZ8tSfz6dHaM2txhe9viPS2gP
HiQ2Tqkm3W0wrJgsf6kqD5reg3F+KcrqTiq1bFoRC1P+pgboFvEZ6scyjHe7NXIfEZmB+SmtJmNZ
Cl+wCUTm6hfoH/kUuOz7KDzVGEsrd2EcSCTTRO0S8urnDk+Mh21Tv4KSLt80VwUtFJcnVJH6ykxf
JOvgZEPaO2GMhnUgfFeLgq1gmoc/yqPuwNJbx8UMbBpnZw8aCap2YqLUW6McvRHHtirMKlstapWO
oE1KIZqemtRrUzUVGfF+2X4mzBtaTSLvb7pqUTCOIcBwSy5X1dQe6tt5XKSAVYslbETI4edByV0N
HRQHtUVirc4RQd3NGgDNJ/ngWB1ffjBjfsAsp3hZuvNeXzbLt8j+TYLu5pLEvZ0vAjS9G5rYUmdH
O1n9apopuh/IXabstDxMD2Y4f3kMWiLCG6tvMBTvt3CNFE1J7sn+UMaWuXNA249NYoGTrc5EklDH
QetyoWmqRfttWkHL5TxBiUnx3PX34ku1dY1WIdDtwpaurzlIAKrsHqIaPbL6lVDY7q0PQxAN01PD
7XCOjwNnfZ6egLVVOk7A/Oc6FK/T11q4vAEnPgKUSlHuwp5rAMht9l2txxEU9CGOxdC/yyqXGHex
ARcYXmTyYhugkbzTglxWs7PGu2oqWQWyUyWPpAYZ2aStviGW5u6hasQYrUgSLNmx+IIm8Z87qfvy
pk41+3KTSrBzCUFUvtQnSQFV26S+hUSqteMXGax6W8zYzXw8fo0/mYSlmvnyM5C8QMmMblzMSRSe
U2CujY0kza4/3SdX22NNCiQ+NzjEfu7ZNJ9e2Ln47xAZgBr+DkVxN/26fcDqwApOYfYcbbvMzeyJ
72K38dFnUikB8sFkUnpndTg0fvyVjqnt6JP16gmXf92cYQNubkKmsj7uazRvuNTtMNJNzMBtfcui
Ibw6rIyDZ5NrhBQCOWBxRt2MsuCrSjj3WlnsbRoLElm6opOVgX4DxsIkpEIbjV9WeB7m7GPvotb0
fJ+yUtAJ7CmlMubdUxug38SppIDAXk+NHINaW1GNrIerwp+jFpmHse1yeEQlpZ2sHqSYtGHQ0Hea
9vngXozd3NFncbBmlLWpwxxONqr41wLEmpYa2M772CGNp4+WJtxkLaaVBymBJY54V2pPCOKs/+KV
HqIwExDgA/8fKeXsX8awN1WBvxO86WTnWIG1A4jt+i/0gQUdtn5eHVG1/SX1LPGcUxwtJWj3xpp1
jUV6To9PJiIAfMfEfVUrpQE55SnNBzJ0fIaZMUOA667Qav+UYbEVRTwHkWQn3EQS3HZek1iRZ5lM
4d0dTRUdObM1Y5V9hO2D22Hqzzi1EWy4MNuf3SRfcsy9NaFAmFyoSBMUQYDwP1MIQB2xwZY1STWC
zHE1/2Urwe9y4d5nqeuuEgYVrlvNJUK7TKsTosd4/DKaVIIJ27Md6OQb4LLwszkHrr7L2xrT/375
/A1SP47xQklCQmujsQIvgsaxTXGFbz165TybCIKC2EhozRN9N65SLCGkttv8ql13We0MaOdXmyAq
mEldYRbeHCUKcAChtPT8H0ZUuHZJvlmaY48lRLsPq1ajRY25diDpDgX0KQNCww/kZOrSfRRuRfp0
wPi9XQVzRsbd0DJndxToCQ/nSvYLEF5uqvuScWq5G058ccWEcTroVX1OkYCa9/og6ggOZEwsIlOp
JBfLJzFH/qWhyzJGYk5NKlxdBAqlbIk9PG8RqpgDYdcVIDXeiuLyWgAwYGS+G79RJfF30QOU8vY9
FeYUokAkFlS8A5QF92YkjE/qixxBkMNYLUWXxH7gRk/DKKzAMD63YxDPrCG22jUucA/u2NiEz4z8
Zi9vHsa6f5ZEKTEGmIaL2I8Ajr+8emORvT8T8ZI9QNoCd/D/q/mUOpxPEZe5pvLCLOdi+dYr6OYU
RkKnyqf0EtFFoTQFiG9wp3g3gjgi7yLq9MCHzZPNHBytLPc3tNZXFohATdnHBvE/sUyjIBrng615
37D/Iry0DrxVH5ej9qweQKrjdU2X6c1I1is91YTWyFADyJJpCxE9LAkJ2nVkxTUG4Z2HQkOYT+Ll
besZWtrTh+oz2t8UFx/+CLRKJpnS8CKVyotneaCJKA0cRVW3VVscK5KAsF7EY9MVFV2GELx/Mkfy
2V0UlT1UXIT3BboQudKzUx2lOJAV1mdUzBgMWV+DJtLntY+ZQr4IeHJL+VshapHEmeemWHOxcoVg
n9pxELPXPOekVQpfe3yC4SCpmkJzcl9+T3VmjfNcWvs1n8jNQyCVX+Te2Q6pjQRBefcuKW4NI9yx
3LfCUYWxind7KwoCRDvwJlGXCRxiGB4XxTsWwMsqBOwACZA2ozyxF/wImoK5oDE+8rpHRXFtoHSg
Mc/qVP6qDmi2L66Agq5dj96I7ybzMMxf6Bww0cd8AH27vu83we5sEiuK65nk29q4bvqHMqPyyoBQ
zBuvhjRhC/CaX2Kkiiw8EpNwWVOf0ur8Du4mbmcEWGhLTHDq3QXKJvWiVZ6p2kf7VIjeOHB0oirE
7xDWs4s0iY2nXetugubI9PlpjqKFXgHOtdJdWSj6oIQdMemrWW8hSFEtiBh75AbIOPQoIQ3dEWcx
sUPaIPnvab8DQWDJ6DNLjaUljIy6GdIX7e34ct224g1Z++L59DIBTqn5ZscJRx0yWxl50hrzAe2i
Ly0hk2VW6xYdtI2/6aHYmZoW7aCrnA9LkaqlAdHsF3/HtMAeXvO4LLvk4FCUwJQwhPfN1jXn4LMN
HMvSwDu8Nn3CxHQARSoNGqeZyhjkn23zjxSxFNjxcNMTCjtco0LoMJ3mrSsUGy66glbSoGZnx+Bp
4RidZGHuw14zkjV8vIKWh/3sakv3ehlcUQU5Ttce6nQrkOXUVbBmDSc+mRIPSUQ//mYPruVcoK+I
KTQ+3wKolSxoT40/L1D37rLuxQnLautC9+eoGb3FmqE7TCcoB2VvRPJbDWjmazv1gYlO+mzWw9eO
yn/1gEUu8K2CxFqcuaEM921C3WLhQ28XJeq8VNF242QRhBEOJcShwW5EK4RV7/jNx+a0R19FO206
PuEBjcgt3x2qRpb9e3+pPtBNFG8R15oF+me226KNsN/M8E6c1FQkz7g+l1qG5mVinbavnXd5pHmT
Z7sytUBDzU/CUKpw4CLvLATs89uO5e0qO6ZKXN+j0RqgWX2lbxu9EGqSLxOWBjGzH8nXX4/OqIpb
dFRHaCdQ6Ol9v87Q52FxqHkDlAl1w6Obv0/PCLQ4u50PLfixKZzorGwhbHzMFrRE6k2Y1+SFGuRS
0OPlmiDuc4q0flS75E+0JlTQReQMM0jSFwRM5/rF8QcrSMrBMgyBAh6tP066S7YmrC2XNomqN4dN
5u51qMSYtmCwYPEslvAnsAdiHu/dZiAvOWUH8NztW0EnuoTFNNG4nQ5nxELdeIpL3xqIuQGjjViv
v12W+hmA6x5XM/Muinnfa3zyGOAbQ3PDphq4BnVkASYqv1VL2Irj7iKcb0wEVEORci1jW8FJYhuO
RTiEQUSTh5wX9K1PO9sYLzwI8/qRRZjlto7MtWRel63N9b3mW1jN9ZCI1MULs24VAqxMGPdoSCiL
P4NjzJ+hGtGkV07SSHlO0pjHizF/5rdCiwiJyR2FRyu6NCQDGrz1NyofwH0jxIFI58NPv5yCwg7m
xWDKfaavbns5t3OZmJQnkqidW6kvMnfjE1pMn5ezlE//6Y4hCwc3Rb4BZu+v7sdRjIUl3R1HvlL3
tEAv0XHyOHEBJCHjlshcVRGDVNxobBxmjNJ2NDl75ZeEV84/BrlW3FdqBgqVOA7J0g1RXLw2hynw
H7ZnB16YNAfoF6jt9QvrPVXBdWGBu7x+lrui1Kys1j2m9JjRnKNbsWFIhgomO06KFWbny43wF//M
L8TzDHdXPUJDxyd4XhEA57nz001V4jgEP3i1YDFVV33ZpErPT2rOCg3QlsEiaQZFAIRRGQ7pB/ZU
esI1xqUV7TlxNkdQFYV78vDor+H92oBQH/i6ZEF/lNhYPmDsFwX8+UCKIiaanS80tMisG+Jzujaf
ZVY5ZhNG1U6FKmfZg8ARxRxbl4zjSkZMDawIuacxQVN1l6Yw6p3e0LbBRSJA2ncwyTfQrq14l2k6
7IFHG+KcjEs/O5nV8wVfECjSsMWDPlhfZ7O8GTB2ktaePOvzJfT6+OrLsg7P9EjEhTgTrmkyMCmh
ykv5hnd0UekJ4BWg4ZnymkgidqAYLMSZ7tKAPQ1tvEUwb5ZO5z+ClI27GoHUx6+n4bflxB7V5Mvl
QccN8RAirT8wymSAd6m1frOHwIqDnH47C+CcrEQkfUGLOyAkeY4eYAgQl6zwORdbsFhgvQ/rC50F
JjOFx1o8LMk8DRYTfJCnYqlyfqDzngf/jZHGDbCbKt7F4UMJw2sUyLZU2AotW4+izI2BUGoIytRg
QibrgwWfDwJAwRiRZ6AlVz3gCPwlyUH2/nbCC//r1H9mxUjMwEuEEqnXwLvE2/03P78LSdCSWTx8
Ifss+TjW2PQEOg9Qe4ioIrnCwAuSFgXwJR+cpMIrkAqyNA+wjmkqVSPAQIOMDHG2seKZamIv7RuV
Fc38YgCEaUR2+/gjqZnhlnesHZnQa+EnCpZuTWopW0sC7A1Elam86gus/GkCCOUtSDpjmmJtp0O0
e7knsVHbEhcnUNkjBOMTfWEP8Q9PUEKByx7BI6fjWWqhalmg7pfSyJhH/CL5GgBbgh31w30j5K3Q
jiq8fvQ+WjV+zD/m9qg1hpeb/BTWgtBtauSrfoNLO24QA9G8CjxYmAHRjT1H6GhuFSgoF1O/ygHK
dKlzKZ+cdzNSQrTL2/OWppohwpT6py9rZxaPodPT8AFur9ohMpbDVF8urmHFgbxMLQCNOTkEIFF0
B5xWgayknSqMWp6cHDtXfl119h5BpSlX8qhOfg/hHpQVIQMzmemqISza/3hQJndR25Od4Yn/txNh
9YWXrxbaGJXNFpbgFviYyUGRvuEwBM4+5+HYM7MwlAJpPRF0M3vpN/Tfzo3J8iqXFtVSihGh8j7k
StQS/65lLKRl5b+IQvS9B9hgtDw7ht2oP6x6w7sRLWht58FVmHiiOtObWgS27r5QoAvxA86cKIZm
nzNRsIdTGzcEJ3gzyAc9JoEzGfH6l7Qr1GC4BCxntxpgpu7Ytf2PJPYTfD43wNeN7M8kA4VX/L6B
xBvrMhH/hRyGoWsvE2nSvHQD4mu4gxcNtyXSJgaVJk/SspMQUx01Woh7547HDri1n/i2uYtaKzc1
461KErUF1dGXR7zM3CMkHi1HgGkfWJB7uHN34S4WEvSF14ZpsJUzDasDEJzQCFO+x7Co2ILfZld0
bD8puP3+aWfwImk07uuDR7R7iUaWj1hB1BdYPhFn5z/uwiQ13EIyWeXrzIPO5irlHkyE6Q1BoItv
0m5eZVrxMoLiKC47juKpXsfzWr6hogIX1svVOxg5uAJWhDUE8QtxNXwTAAC0r/M7SD2Lk6UlN/Kt
Bfl+sgdTitBaLAh/9FHqDmPnem2HN3Woqoh7d9gCioGDHm/iIImS/LUmIdB17KVNXZZdar0VwXJ+
fqv5MPnApB0qCfrBjhHzIyMD/2uMXty4ibQQvVrpkG2sV64KVidHfDioZUaRhc/exOSAbfRzafXh
n1a9CUh5w6sxioMj0fxRRsZ8hwqiHuUaRL78VxsrOr3mLniI4PiZnPNjp8fJNwFNyFOXQplqS2yl
VlyVM9UeaxylhotXAfnxrcT64Qrjmd3VrXLlRLmnTWJiayRxnKkoNZXyOkz7sMcmsEQ9+blhMwmz
HCAVTojJgcatHWYrGhQ1CRkVyoBxwec9KU3MzLOUNoM2XCakNPjjEMUcZcZc9BreiHP7n/ba26zh
kZGvlyS3W8w64yqW/dfAh2NxoFrlCJDzN0HKkMqM8GT6iJ1tvHIEaqG34t31uT0D6WaZJN8x/glZ
uPzrpp5Xx69pb+Ub5ocPETvpPK9Fxj7Lxttrl4wQgyttaIZVZtc9gd/YiGzgw4goS1Sv7IUw5uiF
JPAhAfxjsG0AX+2gPH+osGkvrDeVs2VjPumalQVofhTlU/OwLbNFypjMI0yxUa/YxoxIr9I6j8gr
vGMIoAPyHgqwyq/F4UOwxk+gxj8Vr0igBrE7m9x3ZN/kak+SWvsqeaFXQAH2EHemOKEOOhRK8/mr
13kEiyPs514oWTO1e5y/7kmer3MWqpP6B6b6PxyurKb03u+OymDAZ+ZtffStyXLIJwjMh6BGgCNM
fFTj7VogST5jxD1dubtw2O8SSonyHNz7e8L9oMMMtVzjRqh6waajmr6cISs/D92Dw6gJJv7FdmkT
2IwEZ+rY16oF/qVXEkkAU+8885qcoS+hDlgf8OpEvbWVkYxx9vOq0oeuraxJcXgmfXoQyX3OAMzS
RDU09Vtkapqe4e8xfCBhkRHFmzg/jJP4mCaiO3mmQflYQuEJ1p9PbQtYFD9sBaLRhNGLIgRrICUL
Qo9C5W/6JSx980isAYKfGxuys4HtxNLrVxyHRFi4XNZNEZrLbBd8XawBJmmv1pmPYIK1om3oC+KV
76dOByNNt7wqwm4LPeyD3hf5vYjONIPlgA7p7jkWmU6Zvan7tBxtFpVgqpL6A0sXSM6V0cIxy0Pu
l4nqiUbhX09W+Wg34QimY0KmAkNgSb/tpa3Sy5V7mAAWX5UGZ5bsjIyUxA/gYNtP+l3rtovMnovz
j3UBO6S+7+MjAHYUbZq5HsM8UYsb24zTJqTJZ8kLIpFHmsmiBhDim27M0bu5l18xqE7I/gKFOY1e
AuvTn0nB9J6ypKbSgB7PjSWC6e8ymZQUvA750Q94aQaaBXhwxqC4Gvy/4bGUa+OlXKihCv+lQw0W
8VExcCFjSwbnu148+tyqk6SsZXW/nm+ruowEg72t4zbN+nIIwQHR7R+LktpO8A+QH5bis7g00zKp
Efr6PTr+gmAQS8TVTrHEKMDQpjCqO1iThLIZXc1bK+cPp6itC7Hw526kXRCzXxX26DynhcLt+Lts
i7DmjJqYle+Smtf07oeuf5aSBRn+1KEAlSTkvWrLenGsgUEV4mgDTi8O9ykOT5KvoiMsywyGEZoN
Ni1lNNAnvSECR8xusmSXNTrDUvxaVtUVCEo7dqDQ9gFURKPFGX5ANQZZzI9Izs2lYpXVG/z8GUDo
RQ/GY3rN4um1/6E2Q0QZ/GEfcU7Y9QAL1sG2Jp7tvqPfVzKy4NL2aRLIlKJZHD+/cj+DnXt5q9ya
AnNo5J8bQ0b8Ukj4uQbGHV/HoLnfbTI9bTzQsqSG+f1/bHiiiIEtpMAzL8dGDgHzYMC2tV8CHITD
eZdT5rW5/LVI112FbCD5s/xwaiY5KCsH6ZQZSqYXGVnn+reZVOXeZj5UsgbVodQf15+80HGSe1Z0
YMujf9LXjfFCY7fuzPi9B9yNObGvaNVxDzJhW7btwQNSUCQW8ubvlXc29V8lzaxMWMMYFb1oppJR
WqpguQQ72cB/P7KWUoMjW2HMD3ux3IcXsOgEEcoh1KzYSny5T0oU/j3EWEpVfXtN0NTZDFD90QSa
6YWRXmOgHkS1PvqLs3GKwpo1JqQREBrpDC+ZY9HoHt32OGHTZL3TDc07mvCZeIZ2KCe5IKbm945t
dk6l5ahzsX/JjJ+CXGmi+3qJDXI3PecFCh7bLgQB5yNpSRwUK48H+Bf6QuM5hAUD/MTGHtLOY3ei
Xn7gjC6+rueiXynW9w2k3bZ0ZIEkupdDKTG81gQ9qfzmb5Wbx+WZv5bKg6ZnPyNrAxgRiw4wNkPg
4QFNqOZ9VAKUyT/JGmv1xL0y/2rj9W62zYA7Wm8yve5mPCQy6j7d+JDqACqmvI1HYiICg2dMnJuw
f3PtXAd2HmB2audFoPEd3U2wxy2u4lahUOABaiizuYN1AbchoCMPvnm4lfcCmQX8Dvki+rtSVXAl
KgrxG63a+XfG2zrS52iVTQ2HGv+1JXFEQutK3SR8FqunLS8HvmeaxavyXOR1kM17/G5+yvrkuRWd
kwJ6RViS14BdekvL603/Z23dBaZKr1SRivl7+aiKkg83vjKv5d1rqdXFgHhNXHq4vqxP5yP8F1pL
Go/4SejTjfrSolkkd85yNEJwUQpmBQxk+6Y0C4iqdKo+AYAKJC8EnO1R2iJ59aYGNLtf0iDxquac
UESLiaijdSAis/Hc0MqJXL759//zjrUfaXPCnNebkWUuk7Fa7Y7oJQ7PC8nxeQ/43hB+VNSIBOtL
hu25hAYByVHAYbZ59Tiezfo1OpADvoluTX7uJHX+KpZcWnPKRKYfsARNB7rimKnEcyQ0hltSKog6
YBv+KVBJRiiwFi4vlvcDz3zBLJ2OAulJoDjh4eM+5MCBxJS4qVz3Z2nzzH605GMbRHyx2CAKL+W1
5Nemd67wTxSWkbN0Mkn/PdwSMajGEDz5lwL5B9DbT1qV6bzp6QG1vx4tJ6Jf5jWy+CksRpIw78Te
SVPDAn7Qm5KUlEWu3vXy35F20eritbLQTwkwi575bxzCC1y8aSt4wL0Ztmx6CcszT64P2cv4jUKL
H2NfUl/heFgbcJOXMbEs5mJOl3nNCSi56BWoN6J5Bd1TNAn0/DzCNs0deUQmtUcMlmA45mo6UqdU
ud0qB9szG3qE3aASRku376zwVr+h8Xm1bpzra2lL28cC/IYHOYt55405RS34GP8TeL6Bu+ttimk5
UV4EamYj/QAOcaX7/SYLDJ3ijzYb5omW/ifDkHD3yjxWcNtjF9ggQ43VPW2hfM3yGzvDimsop9mx
zDj/bsJAVqSGDLh09Qe3jd9r/uUL+CTiBeYdq7G4V/0qZ31UEyT5+XNpf+BWvJsV+uN+ZOj4yVgI
AmkjehmhqtgH+yH964sRULIIsxccCRRjBB5f72ijkli6AmaouTvvn2E32QzaFxS6hZjaX0XdGv2r
jrXvQtRvvu/dW5utxQiIgppVowrYZPiF0JscEvS9towcLRCpRouGxftDO0XAdegKr6NaT+wIsuDE
oqnVnC30O5UGr31/6M7O6AK4we54TsH50gUFPgoJBIjQm8yVpDerpSfK+RW9pG/ecYzeDmD2z5nm
NF1OzDqzaO5EeVSxhrJSFQicmaa3ilr45t6UXJCCB0qad+e21b5D2XZRA6bUq3kE4IpIAb3uLMt4
eI1gghjgKlE/F0wov40wq5YijSoAxbXCB3q/LNsSt/xqxEjC54Jxpn0ITCMpTBGbuldgTSPjj12n
wQziWNu78o0aGCZkEbXcuqXUaTq+qRt//SkbCzbSqBN/VMIg70r3CmWW9wAN9jpzfDM2diVYu6Dn
T6lyZAqotTXW2tjNhYpGVUW3D3CXkbFpk11zF1UdBuwSD2Isc58rFSUYJlf41GgBASKgXTQ8cB1f
FMMAQ4oHHdnzehW/OuXBCjP3x3s7SzAeNmVLbEBUwfiF4dwqypswqX8ACBowsGlWXOnReuChvnsb
dVRurV4bjP05hDxVKHS/uYOl1SM4R5EEhJC4kTSxZ7UEIoNAHPbMhnKYHpaITkHjfE0VI4H1bAZp
q+sAD4vbRqtN4AgrC1WyU7IRWM3Ruc/lwlRE3zlTU5/0NzG+p+pJXz+G/U8Xc3nF5Tdw+rpsAjV8
Icb6Bsbuhm4k+wbBeHLQ2tHa870bwSWaUVe8afCAoqEw/eWRD/LAVNWe3IF08hPvkaUCuitc4Ggv
vZPcWbTYj6ml3TUVnbbEYGnn9qE7q/R0UhQjg8w4tDU8pXj5iviNb+jk/94G7WubbJV8ypwHuz5P
y8FALB3PkhRP23NeMWphqEUvOYp0wi1ylMJaF+MTtvuDKHr/tY7TSnb5HNiSvNIJLplKvG7PCVPE
nUuHUH2pn39WQq5ScmMEU4mmhmeCn1PzrYdQQuiDDONP18pXnJOgpHMhAFS16W2WGp8eJ0eNE2MJ
H4UYFTwD+TkHTCY45Bb8/Ys4g2drPFnzxi6Q0cTcLTbWaJMH+/lcghdUxQl8V4IfouMUnik1IVdv
toaux1YvcHi/hZArEMlbFXNo65Fp87euQEKO7vgGimttFVoU8CCHdGIAOj9YkoENV6XX5O0qlfO4
Z25TMsYYycRadicOY2lGVOUYpLEtpugIEUsQAfuF6icWNRJDEyl4LwCV8rGp/bRjFgCwa5GigpuH
fy5EfnNIELXPyRppyU3N2+VqJY7KMyiIq/WrvvkoiJdAJp3we0bn5dK+dYB7N6XGOgaZXzVjdXNE
IWSIHp+IibNOHJle783zWGvEbbY4Y0imx3WjRLaEeaQAJIgKywPVscQkA5VbVbTkoUS3744m9CbE
PhS6DaIQbtvHRuRoTzmJW67LHg6K4ZsNnXL5gsQS3ntvkYHJWMZWjUVlJ/D1/Vh+ZjXxwFBn3i9b
R5XewMfIhYEpC9Mc3DHOTHOwARp5Zdthp44qOP4mrj02qnmX8yDUHrl0u+6Efy+IwINCpi9If3W9
WvbMU/Q3TGcPAFNQ6KN1rpGo1G/lvTqOaE5Qwnu9i630VVu5hMgv6bIwsEznMrV9LR3Dph98esEk
bZ+/hUgPLkIkFwgQ23JIM/EOMAuxWw+7N3UdxVTagFGwAbXu7BUEl+HWViyhKHrmGTe7j8cxtNXy
r1QRKgE5jilDBjpaUX1zH5IaXBzQKVW5Tgf1cVFU+GWXsnHzIfATbJZUE1c4uXpOvjS2zYm5mRlc
bV5ic8DNGnVyl1vvwp0lDlRpqnFPd8klcLe/H2hatQ1E8s3WwE2R7009l6+uxiHV5xshIgoKvU5d
pDlcvBvuRHXnGSsp8UVXhmv8AGtd2otG2t8M4OYeoHOd/eJ0LoLxaH4TdJKZeeua7hRGikKxpXr6
CAnauoskLUdAP0ucypv4u3LiUqIjogvar0bX5LKHOgoHk0NJI458kSfP1vHYYtjEozpe9pM0QyDq
4iv+m80X9E87q2pgR76lE5n8qL7+5TriH/VIPiGwYbwzSUpg+wLMyEo3KkEHsMgNRp9jq6fbzwql
yaHeTA8dutC5sooOkiNHiutaKhSdny8bbfeHRbU9Ho+XkUtKaD6DBP1SfdE9z9S3cDW+rt3EQIY7
ubzq1zO0pQBon/Kpa1s3me1fuR15oJZS4r/PQuQTsGfj3Zt8l9EBc49yMZRNMt3+TBnUPW/tfrDH
vBq4CR5Cbj463DCY4YwZICgn90s+RgIPeIHfAH8UDek2o6DqZ2lipzPBIMzB9v4W2cRQMydQb4FD
aaQvXku+n23dydO8V6i8Ktw9B0PE9hcAyQFV0Hj7KArwrkRe4v8/ALWg7hpn3et0URDtn8HvIgUI
8SkpLNsQaP8Dirvs9DLa6aVIXc0WqFmMcXufc+/J2IMOyfADD2oe3Dx+JKXKxf87TAIK0jCFev80
h0dj1uXRd/BEZ4HgmtfoZNTW/1UEl4ZS5DByDF3utYZPWuCO7YspcbcshpWHAbtA6dXtDaOURv+c
vfDS83Ni/T/83+fy/r0RsU9NyYZgZyfJyfKmPZsDq1MOGbnD9zyOruMRpHA0e0f8Ow4xdu9ZYnVX
IPOftYU+Cuv4ssSKrVLhsIweW4Pw54wo+QqMmMXRoiq236MZT9MkZ74LSfJoN8DuDyUPowzOnCdm
ltYdqsgabTC4Qw9aDaQV61DshKh7gSoPzaD+0b0ILQ4Utndo5XOzAZt36/lI9bvL8z+e+IkAqrFh
tIPwtXWaj38xja/Myq1uL7I8+lELVRdfX+WP4K494X2tB+qB5SDohDfLQYZBpqJTECzFXT3zoHnP
kBRzYuPlGhmEPASFGRfpQeLfw+s48Mcu76QCHbhKMIblPo1j95ANOGLuujTVfb3uRw4CRuHxu790
2yaZiE75VMk9LK2AAz35fZQ/7TPn9zzf9SKvqVcjnJPQ5BpCMsPxdyAwn54+bFml0ba4Q7KdDh3f
Ov8OfROeDEJNqoh6jz76Rg1r/wnwlYcWU/x3AHm/73l+Unqoqrvi9ra/K+qTcBpTAQH47nGwCdKc
/TMT/nDy0ABmFRzuENdjEnLVMhqxBlN8+7MXLtjUm7Cx2+JKKQQLb3X0bWSGERajdA/Y4larykrK
p/+QkwQ7neNf7uY7cKutF73JqSl2JhJeyx/egCI3A6pHdZdXry4TJAcs+CX48SVET4tVZnnr570B
z0sLP3zk6l4S5OuiJfSE1F/6Bm7p0SdTKXxNkKcj7vBqvCw5ZHWfMTFx5hcjCiShnlTmGxXUw3O/
s1pUcYDBLVo4ZVCQ4HnoPPv0s6MZWeAGjKn4QWhzzbR03vJkfwcQPRyZpEWCuFl/PGTe/IM60tkT
TFXJWdCKVMiCbsnmiYZNOdyWI4DjkmZsx7HsesfKYmEKvNJaoEO2jH2ijSCeQp0D5s9cr8sFtYur
Fdx8WMFVhqE6/H+eeC13CnLtvnZoZQjc4XgbNe8x4Dl7pNEF7Fa/TOie259PcYJ+cK9uBy/3Z/JG
TsdRp3BCZ3QGpKkyurfjYAIbT1XwCAn/oMEQ/MpJoKR3R1n7PibpM1NQjcyGdIeLKwrfaO/7OeNI
JpNb/avBGbFErPYMJ3szbv3X44h+f6V23zuDLYt8HjZD0Qu8wLicmT4l/VhqSG0kGUhwyjyp2j6G
cfQ0a6jY//j3U22Gx2/HZoKlMLd6NELEMyggGUnvEvVAN4pNQ68yr16XxrylU8Cy9Yoy4sCTDqfl
AERY69F22BlhuyAwV2gb89TEG1YiFn23ZZ//+PYxzz5PFRyL8TGf55L2vRgxI2KdzaQxL/Fd+jNc
WwKRcaHICAlkI3n4dNc8Qrr54p7iXoKBZf+69l8cwhO0I8a86szf5HeNiBDbT3SJlEbV0r3ACWbP
+4sqNZKr6KxxC5XnYVxHrHqtxp6E6/ZfjiYCI9acZnDSBTMT3Pup4gh7ih9RPmwbGl+yrVA8O2Xh
+tdrBxK8s3AZIN04giVrdatmZwfDziXpPsSFj7Wqn0NEGf/6M4I6+15zt8X76BhPz+Wg9gjVc2UG
n3fV6rKN3mx0atMjPVR19p/rfknIi3/ZnVL+VxCyGBe2jz6YvTMA9x9+Vn2RIiSPRUUAGJM4m2E7
WFAXvF+mJCP4Z42RmprVQ7Mq11cPnm58h4gqZfTsoS6yXELc4KFKvM5LHElLM3I8UzhM8rnazwjk
qt6fFhyyM+K4Sc6FCq4CKizIkogvgrtuci5j8itxpIlR0TGlHtHyPrnCl6Z9OrKIePHWtLB60C52
uJI3BAN8+SsorOzNQtw7LVUF7YUwl/U/0CP6knsFFIwbSzpR+onYl6NoP4eg2yB1OwYv7W5LhAvI
08zpsb4ycOLrqAc84P1MhPi5sCfXzcasCOWCE5k25QNlXAMdDZXyAfoXEb6lUMcSuGApnpSNvdXa
pARMZuIiwHHsL/ym/FyD1tQ57CLOld8DM9cwtUqED4KlIT9hByf/2LAm3U3Z0zSkjN3x93d305dp
BWoey0ShdajF3Fy101s+pBTZQqrmyTxf89YCrl8EVv//R3C9yliCnZQ30P1M+NAJzTtM4zOVwaht
NjeOcBXDp0HyZjMZ/UovGJr4KP263AxRjDeiQGkzSOMDZDavGoEjwQjL7xvGNkn4N8oHLumQcQuq
RDdd5L60IVzWKBvLmqjUhIKWwBWlsamTAe4vfNxurHNVmx0+hSqhNH3DbYPemWLS3EyoZ91/+G1o
lYM2uxI/YZpFgcM2gh6csbvV4jsixiww6GemvH7pCAr3O4DkGph0M23nBGxGMw8FA6FVHAUENH7Y
oVPU72rBRtNJ6T5eEDuVPPSHl8JFstZ9ajxIVWyCypZ0x8sSlwn9P7Qdz1g8f52FeopM57OBjcCk
0plmgHSFwcRq/cvQlMVzsHijklM2Yy4wJxzR7Ul3IIJkg1LZ1bN4pl6e/1rBO/0GatEdqNHvBvDS
plH1sLqCaeLgq3c40QG/RDcjTBcAx6cYPyUDIakj7tEHGP0gSN5JApzzi1D6l58ZruzCQgA3tIpa
IdD3JTvyrpm1/7RVNVL2Q429KSoX4r/orLffO17ISJ6O3iwrWxbSdLbZul4V2f5mpCKkiRnPtaRt
HKvRiPMHyurwajuN3ibWYrdTKEGvFCfX5pNgbuK92V4NOImgYuqmZ7UjoTDHfkUXNi21YCbO1UmO
JhrvcWal592ukbIEsv0iHtptvHI3uk4dW17b+AcbR40J/xaT1tVOvLmpthlESZnZsziJ7tsANyK8
wC1KlxIQykgt2czbqwAJfn/TKFB/P3E3kjfJCZWkbEMbqj+lOG1W9tMnW2ilFl78uYZaoQHdX/2H
LRColh3QFX2ptCpZQ08sCgGZaf2OEVJ8OqLuVjq2PDI+nnuZ/OUHPqGEuudN4+x1RrfLmN/YuySJ
ty4TVtj+5gND2S56vAhWImQA0FFkMASyBxPDit8L4+xrLabE9F1rX2/PfEzqSiXfqzvZlb038C7C
SafJmjXTM0Ea6f8aa0QQj62wuB38SUaX5m2yVr4l401Rlt3q7tsLBXWj13ZA/jWbbjfX3sTBeJNw
E+3P3Yhiq6PrmMZL3UBeT9LF1+0Ie9QfhNWT1H+7L5ig/of+4j/crZ0Yw5BfbgLGAQzplAd+6Zc2
IB5k80Au0FezG9KSkMgqI3d+Vt3qeUikrfFdavjAxBw35pLGwzCgSCcic4fQKRpuUOOKcoEXHbRa
rMZ3qL6gUgrDesL6IjWZTfS8YkcYDFCq/5iESdZp2YXzaThkgXZLjx4mipaE0CaFNf7sTBZnKWLQ
rn88CH15sjvDcpw7zthNBXK4+1hOgeoHl8B5kJuAetvL8W2v52YBL+gfuHgbVajsV0JrXyyPEhcq
MAhVuWwgR91ydxv9VH6nYCPEhmWqn4/xsW1IBLl+oX/WhIfhJp2y5jN7s/oJr5FdxALF0EhY2phh
i9M/iguGj6FpKW+U5R6WPdPjew2Zr5LGI/JrufgZRtlMfAQnm409CchCAu/9B//FKWYBVhnrQpus
LVyyEq7Vnxuw3L+IVb9Lo6Ec61qfNkiQhFFlfttHtEHvaOcPhoDkLqXILbNN8ujentcVP8skBgdW
iN2Pr8nzQd/Xn+xaviX/g4493evKMbLFwQRY8sGX5ewYEe3kdZdhPJgrRZ0OT0JUPPC4zqtClv7O
rGXGAL9csLKrcMC3i0/BKT3I3bHYbNW7cIURJaHDHyQowHWW3YfJ85EckYzkDrR+gQnoVhZsYkI9
dWQV4nRIQCVcW9HzSRoQBe0wmckRJWv4Pa5zuJeTjf5YqHAflEoIPmbzyOFejzGxT3bb+l1I4zHd
3L9IWSQVmf7nyl4LswOPFwvidh4UMIsGIUByqVydSER/jqygpfXXjtGPcWXFh3z4V6GYsc9khhs9
6B1GhBL64NYYce2r6w8/pKnQy5opwRIsOUJv3i70ioaLrqfPpCSnLyxnJapODzRtB7Gd39m68P46
5Ek/HVvt+QcZVmG0IOqJraHeOx13k1prY9BjOyr2XY+mFrrdyLJ017zBDj7DBvRyXA8CYVQHk1gG
GyrVbjY0XFNlXF+938DA0+PzQf5WD9GUScdJOHXgRX1065/DEohtFBJ6C5yKY+h9jsEKfRaIFB6E
Z+3o7SMD727hRw66YvQp6lDFXI8HwmXOl8r+gRQM9zdy5sQ/4kueNQP8LJIUuBmIGOMaeN6BZP2G
PO3e9MUA0+NAAQuUd2lOZxl8Y3S7tU/ShZDT5sLsawrd8peeCvJyRNL5v07dy9uLSMGqUR7UmflC
3ymFkBoVcDm4x2HK4LzX63pjOdP4IVSfrXwMjJUCckMAnYmZT3F819/40TG6Pb46fPsruf4W17l2
SNlRS9oTboZmBDnXBOEOsBFjs2kGNYGbebEFi0PJExGNzJ+xe/TPOOtfpD0fc7w018aOvQEOtxoQ
l7N9fGivZ+U2xHs370ttbhSHEU+Ncrpk60gLYbG4lMjEhVshKKZXy4YDkOOOH41o1f6n6O1AYAr4
mrcxyzCRUXuM6mX6PvKsl7dUIoJrrLNxmtJZryEq6/6NKFiq6ADToSCR8RNWyUZ3+HOfa6gh/UYP
z1jG1MkIKozu41m52Y31TywqI31h+lMvQ0GCuePieSqS9boBKA5QehZGYDB7/ayZ8PKFDZ8oAk/R
IVny2ehHmlFVB3OqD93ChjCuT9o2v3/C7mUWeddHutnqd6LkIIAHn1NfY47Gn5qWPjtJSefZRZIG
/v4z+EtEsK6wNFmJZWaNcddNUnQ62SIgxevzt1zVOy+eer+Ekgjo1xdDBeGVgT4Xc3KdDMwotq8P
1qs0UuqF/d+MeWJCZ/EG54Nj5wNn0F8z7hDRjVAUqIcWsc2WfkftVwfmP/mY2RbplPJMMsgyqaaK
hP6AaQ/bjAiZKSCpl9SYr7eAyREwoK9Wtg/yjZFxJVHyK308hNc4xN2jnTSZ5IdkpN7Ctend5idW
YnE4XCeJ8W4uPu2nLIv+bo6N9BI6cQA6O/SLYwCIZ1RpZvv7Q9xN3Y/Fjelr0xQq5gpL7981jcvR
MeXlm0uE+KhOueMWgX9/RvudMjcydcxjMZPjlgR10AYp7okGQ3XAIOizoj2TWRK7auXU9zl9IcvT
/UL4hIa3F4qKb3QQX75btte9JaMEyGaUbTqQaoqWPcz3qLbXSAMGwgog7H2SHw112oUElTXmhLEZ
DUO3smmwTvuwrib3HVXRARp4BLYlMPoQC4sjr5A8ZuJuI8qStOYAyIg3M+0CGb15mb9SGdMjOJ2B
ghtboEwhETQmdOSE+aX9AJjAEkeofvUrj0idA5c32O++klI2gUXdwnrMgxtUShTGGz4SYDliWFeI
A2E69gKaEZnDwHrUSOMDyh1t7CkPFjSTZK6TW3TcHB6lBcBB7LI9+nXmbMzZfSAmcpYhfGxjU65y
SuLi8UyH7+/CcVmibaezLVj3uixEYNCF7l76ApW4VKL/jGr0Xzh3jc0qP/c/8ihtaxx7e8PL520o
jbRmd9Wv+MiXyA9JFm/TFtPUGppLLPGThIIMJq9J29I8L8nHAtR6xnIquL/qhsNRZQd0+GwwHVJH
fZLqLphFl2uOrjHqW43mCK+s5M12FeQwFrZf/Ewa8IK/yVA/rabpC1JwDF9Qt5vecRJpch5WkmXj
VAc8j5JOGEcrWAirb3N/eA8Kd7qB1D8yHiqeSCUbZtdfrW42wH6zrFiI3kD3tMos55HsLew5o3x4
aoAFNVb2Q0XGqnLjxyo8NovPuRTNiQCYdLNzZ8UeqyDBmxxapP/zZnJm86bgQm3i5KUe98SsQYft
zFcthI3REz3qz58LOYWrES+6EiEn6w9gXhUe4CJUVdz90DoG5NrSkQqYXS7jboxq8gd3q0iZ4VFO
ujXTMonRD6A4wcz22+Iyc8HST+UXUBaswb8gARbvQaALLl8FxFFuReOfQXRGhrutxDrVoKkTqkBg
lB3ogmDLnnFMg4mkMmdAYzIXzHPSrrh8JUZjDg9k84kSts9ufS+5BSj1RAFEghYERDzJCaXiyV2h
VFjN7Qs8tQ1v4T2EvYwxyjwwUGJCpHTz3VrUN6lXSII5/hkS4kXIZkn0oJ2mY7eqaMMKyb+p7xvC
68fSyCcTpGtbEtUhin/IeshR824kfvuryktCwKVqQOSPz+TM9IEF9dp+UOrrhJ31UMTPuRZ1i9RN
Rdy2Nmyqk0SPFIeO0xqQJK5xEGc0STVD4SxdPeWd0vVCrD3cQ6R9JmO0fbkPKVEpgKW7p7QcK2OL
hvGYdqEP6G5lONkpOmLbkeS5eaWewyTXneGFUfhx3Xva3o82Zx4c1cFP4gXy2e2uj66mng5Mab+N
2TZPF1tZ3hnEKC37c+EbWAYrcDOtSdaFaVqkcZF4A7EaLHtS6gkxFY5fD6MBrdIPNoBRpYdDpxlK
uckC5b1Tvi+g1WspQyA018/SjihHL1QasmPnS2i0pCYklNLboIylz5bSZVYmgGl0HqvrMoMB2VMg
p3XkUHfMGAqIHk3rTH5pqitZBF+i6X3RTuSYnvpSZj84XsC0kFd+XkB3Q1DdjLCm3rhnqNQOsdbp
mKHTRYyRwJnnOqBUpzIlpLdD9LpFZavZVZOUgOo35e7PVgQHixNvZPvX+9EH5pW8ni70zhxalRkp
axoHjslvkuuWOT1f/BEAT/J817dnQ1ZrsFRQAzP8RfJsL8937ahkAErLxlUEdAXwQryiBfjkFVtM
jjvH6emuGNTHU5ROIHsfzTLPtKX7CL/liTzFgTihmNKIQx1bw3XZcc2V9qW9xqdXdsQtPWGEU+HB
8Q+HKa71uOvb7iuIw+mFK9h+ENROqaJESQCJO2kzMRrzELmZAepSIbFr2JVT+Hu2OygzrJYMhiMu
b70sFgZBZk2w52HQd1SGeDyVlv0hy00N1lfP00lcwfCdxDPCHdCuldsj4zdNpSt1G8mKWmAju0fC
5lzLng8zKEnTgD818mXD5tZSY03iFu3/tOajKgV9MbrF+P/FFP2boE/rI4Fs92hF/b4kbKcwEEQA
2pvpj4+EO5SHzVckQPfK5W53pz3HdNNHXB0snN68ltKvuSZdxA+gg670WcJs2WBVaphYTGu4xT3B
rnAbjp2eNHfmQWgbGiSWacpsj2dcnoVR011UN75gVNNqq2ItlITtvLzhEXQYMNP5dQ6iCfrumoT5
tk51qCpuiZh8izpku7ZXf0wc0R2MQfOQyS1/BcCy7/faAqYMBCpql3yfrJno0fgAmVbCe8wI13xl
26dEWAs49t/gGOm2tKILFWy7/pPpVZDbP68fnONpPhNxJhORo+P6jEifO4F/UwLEssbxAcAwq6xx
u/jw/QW3FDtrXslSSJy4FbP8ObMJXAFwWTJiGy+ibEvlBXgxmgUL0mvv8lzdwdqIQBoVESzgq9Ai
MYVj6WMGIdLGUDIIyzxbfIe2w50wf4v4gk3ZdaGjKWalAFv1oRBzzYTCNItnczBdJQusZJuSvTc2
U5eWkZQlH6ijsQrAJmL+Grp55QQnbe2+jrWW71Z7yk6xq5FrIijZZjlXWGw/dKTFBEwDR3RK0R/x
K4nJttp1Hl7u+jZRg+usttfowRQdq3o/Hnv0lRGUPIkY37LIhwgxszI7KQ5xTqgj2qoEMs4Sf1vN
/5RrNsM805pLsbW745Kt8fzmey3vaCJshsb3CwG/3BZ+8UQNyKrBYbFPpw5kWToebLSyGjfJkHUL
84vX/9OsFL2+cjWlS3XyMFAV0/bSifLuIlaPjvK0/UlM2MJF5YxWBiSLRFVtlhB2t2/zrwKHTfzd
Ea74D3sXftBgAaY7Pn0n1APbVn5rBC9YQlpOs/HLaDl900xg38r+m/8Dv6H7oLUvVgX/Wa6dxXsV
J2jWPSDzwEoQNmoZy8+rJq4DJFiWKx/5kmOHx7IjuX42WQpYLqBvwA3Vd6WW+wYzIk5stWUYmcH4
ggeOgrQdE//dVzz0IUgxTk2LywkVaQfv2X7Q/9SkjlU9c60MgkP9TLp3/7UPnvi8kV2J/4Fmm3mU
NSBit0Rr1Sl4kfx0Yq35QV9yWzIppjeVfgu5+kmsjoiUKDUYpGWy3p0mo6LnxtpZfwX4UuwCmRMF
Zifeg4YHbxTTmkvy6RrR7VY+824HCWKF2jnm1uWj31Shavx9wcps7XLthk11LEoQgQd/IFR7U8A3
hhGumiv/1f3OhhxpLwVqJ5thJOYFhayMkB1USvb3SiQG5hyXBcwSL8Je6hqJdslV7tqfRSssy35w
DRTZDd/jNI0Yrh/EQgil7Vb8bunoYgQ5/o0Y6oBYbcrY5YddiehcvYLTkmEPRTRsMue3L7vtwYUW
QWdCW14FHUD/7vv4h5K3S8YHjmFYRBcmwIONFzrgM3ZbR0PaBSCiNj7TMYDiFHIPWpz4szcxkqm6
+I83L5b9JYdTXV67TmZ5SkFyWI8pBF8RvVwsqtBMOeSRkHXNeg1mxzjUQl1BZweZZzwszxQrUpfF
lmdgCkX5O02tGxnYFdpizSUFQCVK9Bv4utbZgRaaEXhvGanXVGB7VrcSHRM3RSEHeCWqyt/jhynS
aIZPR7h4s7xmqUgbuCNny6wXbKt/E+A2vbl7q3kyAYUWyPR74KGw94W6lVuE91S9BW5dmiZbMMYT
TaKnrHlGAkMfimJ00dI8BZLKOpnMFvF+n5XbuBE+etJWMfFra4EbjUbdo5gzUWsGdbO8WZkPRSIs
Dir1F4fPRP5qSDZBxTIRDQCGa1uXxcNXiXJgFRQecWmsAOG9sjt55ryAL/prC3nGRyPgwCDKrkkH
QfiHHpp5aL6fgXlNss8NYN50cFXPB1v+LThKzL9hn/SmjH0r9bo23W3pdLKLfFQg3wEozaoY5i+2
OlmjnoBfIfl8dJI/cg07QSlkjKbi3h3gocbTvTxi7X4u7AnnAjKJcyFXW8WoONPfnByMgKJ8749W
IzCkC9q+wynvo0rlPFJvVF21DmNTY5g1mS1HDZ0EJ7OzGMMBc5e8bjb877XOiAdRzT93riWOISDI
zpcp+ao4u0Z288iH+4w69KrnkpLf7bDHe1jg9Daqb9B+BEB2RMhGwkB+Bidw+qKb/xC1tluQIrHk
8bXcgH7Q+HRi2IUmyB+FStTBaHtX7/Z4QVlNaJqk7QJolBR3rOnqsSsVpUTSkrz5zPBd58Ac/pEN
wR+Kkh94CHEyoi2w5fAH+k96sacfUMGhRDkbBJVX0/lpTOaTTYnbvSR/i65uWVurnAPEs490ohIO
49r29hEk2oo5wYlAIDur99bNgvAkJKe2b6dYuKXIdwskc3CVQ8hs7B7chAlnlpK8s8owEZwibzpb
TkyN6CrmGHou0d3o8Gaf6TyzyLZjXkmQ46L7kOlhXe8aeD/hR5cY8g9nkHT4l9woDZac11Zcv9ri
Nuaft8pfXD1KxYz9Wrz5b7uf173I1EsHIzAjArhvpRcnD6/vCWqNelxzndHvI++Ro8QIDSBCqfEv
6Y91NBKy5jEywECs6fEhvWYYSCIZL72wx0WC9YAJXB77CQEdL2Y9UfVsZQeC5rupi4w4H9bu8i57
5ThQzbZ/lbfGfiazmrVghortvZuFjXzylElSqOVje/1cshkox8jsmBSq9rHx/6HZfGlvOX+ckpYD
W5UfoTmZ8vxivhxWlSEYa5CnAmvTkpHezMYBZH+IFHRPbuT9CBIhqG8HN0pQeKsmMJHviYnlMWni
TpsSZGRA9S2jV7iP6YTHNYrKVGjsHcXraIlPGskF6gvywt+GHry+OUJ+8xKjXcFWsWiXi42ubCGX
RhnwkXsfdwF70JTtgpYrV3etM3FXtLgtc0Y8gxSp5FbopvD71T6wsY9TCgrQwuqPotZo82mV947E
Yjq/SpZgQcOtvGFO0omqUoJjR2HA45a5wzCaizfBofbJ4mRO3yh4T7oc6XSk4HVebULajub2Rrm9
cSi5pBCdzyQ2SprjlIS5/tvI4nH54mj04DVhRSm//z0uVz1M4iDKdswfpVbPdm7SK6Z+mtRWmVVu
dTPwnNZUtdF3sPgRIbS6SSSmBO3K/ejGLDPWpxuBhgO2yymOWTA5ekG4OyzEobRaMgJ9LZSDirVb
npHId0FC8zCuumSfWb0vtClgOVJ2WmEDY3+cmEyNmP0bIgqmSy7wreRIZ+fRrlH4PuUEQrLLujjJ
tJ+RWE074V5dhWbw1G9ME5nmwGUihGYI+G5Eux+qoGAHWU/Rb1YqDc6DyWRbWZlbGFj7YuqGCNYx
GYsYqflHmAexgnqgK6md1ZxqPvjMpCk1KyFA4S3/jd0acP1+1esNaO+Xmm48FVqP3AT7X0Dk3pSp
7f6UWzxk0y+cXGxQ0oNY5BtAWENvz5v0RY3jvel9l1I0ws6q8kxZ9ngemQnOaUDQKJq1GV0SyzUr
NvA4oQEeHtKcrD4ELSJqmK1UzaTEedXi7Ci7AqGyO8NNzavBhJmcCwTyiWOieXNe8dubwc7cmPqa
mywANjTODJqvlt+DqNdpe9aYBeSCm+l+vHm0XIna+YbZJ3lHWU+jN5dUbYB9xyuuckIhRyZa9/58
WYWcLj7mSpCGWaH3YpDMTcsHUqAKwyQ361w1fpJQGTxVVldTm8ZZV+BqUFzovd7HoHwLs4z0FTyx
VvL7dz38IImk86wpwrPNvxw9QYQcym5rl6dWojGr5k8hu1mnV4TfHlEAtUXfBUH5rbleXRMdiquC
kQuRcfnVJhdvujaTHFv3kf1FvsJg3fx/GpRJG/ac16nQG1o9uSUPgt75gZ2WYhkXSsTmF/d3cfCu
QtdhvsEgkxLF17d3RxhJAmYB5pkyAKLTsLaSOgxdrd3bhFCasm/uc1M8NlPjjwR17FrkRusGg1KZ
sIDvI0FI39w4yhob9/12LzxDnJ5Rrn8WeUnTVJUKXRlbfCugMvOdeYjTbOXbMYi1aDo1J0WnS4RF
4P73jMqpE/QP3r+ElT4xJdQThvaPFJa7TiysuQh4hk/RkcIfJa7qB2vdVSFzVe4kUH4nI/168M/7
DPx1WVcMuKdWTdRSfF7in2/Ec334vpsyCPnW8cVFSRd5Ygv7ZtbSGkS3Y/2suk4Jf7rsa1XzD0FL
f0Fy7s6v9K/SVDk6liNy+MmBL66miGHPyIqGDSp01gdq2EVyNzTMm+QU9ixMwHmv/LD7HzRCa32g
X/LDNNRI8hXPt32SKx9kyViS9/ADhkoHYVlen8ooBMuoQUT7Ebe3BpCb+JsJ17CQyQi4g2f3Iltn
dF1vfDJ8Xq041hM1O1AcQ1mVTNTSMlnoNNDRDmIdymTcH5tW15PsAn/0yp6BzZrH/5TQTdj3TBff
2QEAhFAEXqEsmfL2XjBv4YFJpKby6xZ16lhyesao40+iHMHNgZkcYczGuQ5sgnQCb3aCXxTshp1Y
dcgupBkZwEr90YfesXSg2RTlngjq1CirQAV1yjcKkiUL9HjjdHzree5+j002iTR1C5TD3F9dmIq7
o/UKnayRm2MUONgKU4xhtGkDMsgwAIQhFvGgjfyrY700EzaHk8m/wTu1xKYFK687jgeJY+ur13Qz
QPeklenX6CUJFmap/WiVvG0JHDUe0iN7WgUcvbfIMz9VCv/S8i+7OTzoApw5Y9Q80R9RYN8ckaIV
6UNCWOtP+ZCYwXbAERQo/hEfmBFQrh+ggGCnTQlANlrda6/pC8chOGdB8JqwTdaGDNP/aCYW3oOJ
CewjHomPOHfA0Dco7ryXRSay/ZBKIj7Q0h4OZHA6MSVFjqHF6saiYSmzHSaTUXVPNadM1li7/Ah/
oYTqSisDY7pogEP5/uRYE8DnnJAWMlnVbIAvfxY+9GVmTKCOuwp+OnCZLJqB0GZ5edwrYxhEOF4k
XfUzTFx0d2zob/3ypDr6ax5Ru/Maf3I5LLOgC5g9cpdUkf2p3gPGUnD6vzxbbrSXOxiIawOSjZDu
nad23IzSoVjTGbRlo24ibnFrV0dWgC4mMNTqAHz6cPyUFRu09W5QIKTAwK3fKX9ilcw0ONAZvmch
2nAeJAfAT7KxCv50EnequOMffWIeG9qtURCLE3xmqhLm26+f9pydtxfBI1i4/smkB6j1egqNRwi0
n3pH/FIEdYab+H5m+Bh6QbdfaDBAXbLJbHqz+tQ8AAzpsoDjvSmNfsFCsi8haoewTzekjegTGydg
8ELDt/fpkrdZ4x5VTjsAKYkFkLKDXwy4uxIEOJAzxdKHyfaL/cF9Vgf8CkL7/P3g0TxnjRBF212Q
MV9qpUzUuTpGz3HLazV5WIXad/TRg0zTcYCSlqDCOTO220kc9tE/VGAelbV6ao+p2Op/CYfH+xsI
PTRwpyvvWzzNiYkUzTHvdjfUQoHedSIuNS0dSef9vF+JyGbp0wwSgdb5QligGRPDSPzrwj87AMeL
wkgNsb9PY1avEU40ykrfJ4kiVRylbD5PLsOXCfPJEbnDaLz5DaH1YLAewLisRFZtbFeCuMg6g2oU
DPydJRp5QAY07LSVnhehSrwY24CUoUvHf2kt3oNTGS4PjsGwrHQlMHHWEq39i+WRcJD8PE9CEFby
cq88nDjJ/+hhOTyfOOCyR2e/cmYhXh2GzTEXNzboSzKq/Skrm+CdStjImfhvg98a94gkxZkRzAyc
x9kPrJV1cbsKn7+TTMzNGoRaNdjVGqztk0NlI7E5qc1Nt9480ut5TMCg3CS/wUWET2yW6JNcB4sR
9FFrIN+aZhvLQ+tDPkMZbdcxo8IB1Ty2MXBJpmug9XCWaYg0jX8iRDH0AK9emGSDuIhcjPLcp85j
Ro765IPS5Zq/wlHvLwIkyn0HB+E1qxftgmRrbcZQTPcQp1T8+RZPAqhZW7oz4mvcwIwydY/AEO5g
5ypQZwA++hewb0kStPcJRAF4GuU8urKPL9cg1MoVANVWJwm/oyKXXLUVkK74A1dvoFdE7qiI0FzU
Lodz3QQqvrbYOnjfT/I+IEq1Om9T1DU4x0G4UvYwl0NhjjoLQXpE4r4lGHI5ZKoLKfOBHkub4tPu
00pcBF4909V4nSy8D0zYmKtv28QJsXBiD366J2P7IzhNjllcjUyftjBr6kQQ4zdi8XmQTwzJA5Lf
A8nMsOrr62OV4XBvIkCVJtZjdRl8OWHuw8yVM4Dp6SedI0HjH9Cu/A6xku4JLrocEIiAfdhyU8t4
gus2JSN8DAecMKVDTgCKgnisu+8quVtn8rtUl3015dGOLZ23eaqededFrhH7j0o3nxAfZj05y4gO
y4EpYohO48bs7175tTkBP/urOA0FjnMUUayz1ri/gZieDhc5DLy08q1V2qBE2yYHWHU6S63PVjkd
vrbJkAVwISoJY/Ixt3mNXMttpr2m35Pey8uKjkeDa9zUdBHnqy6QBclx8pbwtTgSBJg9ze+ZloGZ
RPMw1nLfoeFJZFslDX+KqmLkL5LA1kmuwes9t+kzedZ0t4swrVcdjY5l/A+No/lYxt/eD90Zr2VV
on/B44FhBMZXQizb8C6UkAcCBzOVzY4fL41jcwZY+xjimEDvrHatynQQOrBKyb72Gq/KeMm4n6z1
IyDCJBNawKefFfOWUV/5u0i4vniEQsmpxdsj23JT62xN4DVleMx3HTT+xERRUmJ3IfgtugHnCUj4
c9pITqedGZTbM0MrhgyOg/a1tOKQOWE4dMm1PyLq3z8VtmmKfG40hXp+V3AEpMD8KkAlricU+kqe
bqYeL/XiHvmPH5yuvdLkUznAy53u104Cv5hLNHKY9QdWTWG1OZ3GtEjf08baXhiSex+0+dzMjJiu
nEh9C4AiI7ZNxlUg0CWD5igktrzixv/qaa/6RoK+qQrp07iU15Bna7fcl/uTdmooTXtFDtUAjNzK
CitTvAbnsuECi+oerzTk2vFMqf6Y9DDkMmWUN5qxyb3e/vaKYIW/eqauFkK+dUiJIpdJRZU35rPF
b9e9uC4gg3dYgbkOp5HYGS0Il0GxHuNH59VnU07F8HXFhUaYLlfc627IsLAp+jc9aSC1btW9e9kC
aTjIlq/4jtOrmX9vhiYSxAD42FrdaGXeMMNQC04mHQEZzwo/uCRRYFr4zLWynpw2rZreB/+JVH2E
PMEPSci+2NYuqhZQ7jdi/MpsXvXKa7P7KF0DE9HzwLPw7vJwuB7Fxj31HdCVtvND2bJK5oQjFmFS
cZToYpkZfHZ/d8KwjGA/sZONRKC/kPiwGsiMmoZa6VH8bWDaJAJv/3afmomf8xTvQRuic9jiH3QI
/6x8o5sCR0bYEfk2KN7DkKMP4VFb5ah1yeWWx6wM4HEA8lQ3avwcYJ2fVxq+edW2DMrFRUmg/7+T
Ua7XxU2gIWmgXEUDXAGC5WSFVqGKLio29j5KM4qTWoZ/0jPG1UIIX+bsBnNSop9xtSfx0G1/vjbV
QJKDCV+qWqnWl8qvNkX2hrSUxNhjzPaZFgU1SRA/NVJEspWfzqFjZyvQYnLw2U0amZ9g4/pAZrmj
swSYJg7sJZGwNVcXZfWF6K8mdBS4KGBFO44HRgLJsJgoTquWoLe5Bh1xw1+AUi+aL9924GX+QrPq
85pORTvfGoUM4GzFqPpW2LzJnkTlH4bbEyq5H8E2P1MZSjJXeC/vY0lIG/CFhzFhyvodYKtGwpaQ
6VCJtkVuCZprV31knj5xBk21HOu9YwGRBMwzbalRQZKdVcbkMumrjxcwZ+OuH3zaUlUWoI1D/s6B
Ul5ETJyt3VEu5zv2ZIMLTpJHH1DS0tXznqhXR2wzrD24pfP7eTf6hbXn7v5EMVbVWsAKtvtP7fez
sYd/I1jd494D3zHBGpl7lZsRmbBZT+xP+g7kazG1ONXLEjOs0GyI+9lG2mMWWkAj/VHcDkuJiwll
z/d1RxQ8K0a/sr79pHOq9WRKOnkFhbe5YegIgYyvR4fEqqkWEHT2xQiObdqaAoVtx5lhZo0Si50G
W4ZrCOZ4d4SfGycVWqMJ8qBrMRYl8G6720I0TQQZLsz0OgJBszM/rknMsjiNQTCH0ss3fLXN1Ybk
lZ1eZoiZTMA4MKqpuFFSJztQ1Xl5Cirg1Qptvpm2R8KPmrldZTLHFb+xt0D5D4Jh/weDC1/oBYXL
Tk5AsSfwfsU7BBoYnZI/uyhFiQoEBSEdnosAMSnettfCs9Ooxtg0PssSLmy+qredQ2PsZ03VkbQi
ZIMWweyZzQS+m0Oz7YO00ZWDy90uEtk1lu99w6svN6e3BMv7yZcG+3G9Bo99KcSHN7QqMenE7WAo
cB8mL9SNulCiC3zOebwgJVD9BSuVabOWPFKzoeBWG21DaNx183CLtKZovAbxPMzd/+9KLE91q3eo
81FLo9rvNGPC9LSsqCqfiLt9zewjr3tD7MQ/jc/+pjXvk/0BylYQN5GUZDbFMKEmH+SPXotBJPoj
3cT9aOIASK7IITJ+czJXZxoN6ytr8CMuS1s4z16fMeWiik12XNBnaMQV7R7uyzTFV8cle5ph1LC+
qY+TdDO65ebfGvvp6Gv+fOhzqSH2LxYTGXzvgG53Rwrd/h5XrNh1vZofwgl9tvTg7Sn6nSUxpC1R
AGQkne1KkXqja6ko5XK/qIkYd5CIQeXjnW4AdtUZMsUWALg6C+UJHUOPtmNTWp2TZVqr2HYqqmy4
iVj+yUKuoc9zJLp4VRwFiOIW6eHf14AczhbGfplooGsBGAQ5ZSaJaeDYebcaeq5eDw3RU7nMOPUS
H+SyDmEYEY6EU4jARpv4YYbVsHSo4d3R4v0e731tOvMTQ3rRTsrOoCmNNopwmyfVRxr4KU4bnO1u
zAOy1cqImlRKcfea2E5YtrsIWjaLkqSVhY7tBFJyfBveS70k2/VueXolwTMfEkoQbAPJil2wY1Tz
ZKcGrEzDTosH/wjseDZwn5BI/YJShsFxdQIsg+eWgwkKYoiDCXXGUtfOMP0fSPYa/3tkUz5ywjBH
TY/Il6ELoOjKOT0lwkn8hOczwMGdRlObeBoaJ3q1f443kDgU+9J5yDSfAIQkOIb38E/0aVYlxiwP
d26HACpeitPoL27kPHDbfI0QITLr404kED5YYPjJDVwqjefTGfmK8tBLP1qUqfg36O+Rv/tfdC15
xQLcDjaaQxo7TRoKE3CuVEdZHbAFaIeJTnjJvZgr43SHKzloe1MF3EfY0QnekVIqB3HbYuAyB42t
u3AyVxlrzp0WIOTzL+Yq25ukXS5X9/kCCzlKEUy0uL1YO/rlfNRhuhzh+I5RzGlYTh6EfhAZ673T
1mv1CNJHaoegezCXosDOxgXBIS1jUIh4ldkf5VmymfLW7frajryGdptNyyfE5pk+B7WiYnMwkUcj
CPo1jzd9gkUt4MwzoNq9x+xhy2ePd7a+5TjUkBH8CqtMJLPMvpP1kjP+uxxtV86hPrxi36RGHkug
mX1mlBoN7D6UaIVGWExDMx4DgEwAnUp9S5XAsAQjSiHrfduMM27LGbt7IoKRxVG0wh2HgMmH5MYu
Q6lZBeSFjjEJYOMogawRseTWlLO1ZBdyP0No3/NQDZUFjviM0r6ZqoOkSj/0/gyUV5BiUIooGDox
gGTi8PhF4RsQQh8XJxCslErylnOJNlCUemhBWy36ZntG/awu+WiiS+cgx/QM4m/rgHQaLf6Ek5F6
dfC1ECAdvJCxf7AsdDimvaSuY42ohEwIwSNOpaJ69faPTAiEHKFq1yGS6vGYq5YOSHDb+TuVZORX
wFK2bVrbG6CneEwePoER6PRwirWT/yGBceDg5tJqnpDoEcsrG2FPkLj/6mUkKiAeQNTzhsUk3jWw
U3QftrRViOAaRaHaKSa4CfC5mBFVzzsHfBKM4CVn+Ha1X08BlIVudvfsRjfTC7BTgxCZ7yRBYTDt
7ubKEqC7iPrtrqllba6NzUhzbDYZzFRi0pvj0YHjdqAKcavHKQ0xre59Xs4abZUbHvaQQgBz5PUi
5DF/9ubk6QiBSm0N9pt+dkhDNa0+P06xemMIjtLH/ZUCWmSP7M05bF8cYNKcyvw6QEyGVpxNOse2
0itSBts2uX+xhE1/Addw8hnShr/T70GyWzNsNXvsH3zodmDCz9aGvhJda2Jp5TBtuX5abxFRgj8q
8WEilZwaM+jOqbaFCMYx2sOZZR9GeKC7NclDs0yv3g8W4U8BDe4oSD13Du8x+bQo2gsdZF4TOhio
sk13Fh4zW16+gr8B+WmwuZsOyMGEp2lGlb/KlzLmjsqq3ph9XjbnF3PIMcUmG3TQnz2EuCo1/eMX
2ngi2Fyxyx0wN2wrBBVg5I4XFaNAZiXF9b82ynO8hfSct2WgJAKd7artMa/5EdTkj8A+W1KxTZy7
CJGPsqtyM50ABD9TCJXbUfO3usu3qwq9VG6H+ttxaufx60SMYsjr+kvLMFILxViy5eOy2MgrvWOV
N7CyLMQtUa1Hw8B/jWmo7Nu2DXAdh4eQY2jPEF5Q6w92XpTVnofNdJG2c36o/ztwWGlXESZgUxFN
wA7b9fOawz75OdTq1Dg6RbQuulASG2vE7Dpsmj43ufkCVw6WesH4ma7hEycFFHOQOtM2KZ88oaoF
T3ZeIIDuGMAVr1VUT71nKfhP5cSrQgRZWHRwtUp+xbOWv/pVXB3BEMpNiQLRAQxnIpWy4N6X4UrS
689SxOy4jBUbMzRCNyQAyR2XIp6NfEfh1M2NKgM/EGKktMRgsRQQZAh1sW4b1k92fdq+ql/1mgbf
eaMWkjCrqWUW5a9lw+sGNtGMRicHYYYfOnVEaPYVr4ew4tKKOR39qT+GDXrCAsAPCClb/DE1CK3C
HemEZFaV1vm9Fpm6nX76yhgp7Jp7qVcMfbpbUICgSA2DaxiKxI4iGnfIwm/4rr8C7fwvUUmcl8ni
det3iTFB6Wm3V2/TRf8tIz037tmINqOi5ZbeHp/5SjVuPUV3NaAoyjtb5LoJ1eSMu7NgAYnDGyxT
qnF0fnh+qtq6WXO0mgYgCdo2Z2k/MIt1E3bTJPVSw79MyGglKr29gAQgveq9bRd2xwQcw3hR7sTC
DhMoubcnghj0FnLdtM83Smrp43tMsi3rCgFnm6WFocQpwAuk9MangDmQdLos46c1HdOwCX7rLJ62
QXBA5nzfw9YPZ4zMt0YvHD8OR0TEES47R1FdHQpnXnS6C8e1WW42+azHZlEvVjwhn5qBO1+t6aMd
G8f6lTEthjUIwlWe6bUqb07Ry1WAOrmT3Nf0Dl5ZJT2Ipe1eGRBdRxlq02cEplf44ObO6wEFfQfC
+XcKpcTJnbc80pXFf9V5VSaD8JGsw8ZVhYncsK483yel6xV67R3HmbMO12zIc4FqUgEzvDsGC1dx
UtKSxuIPPBwI1aEgtEzvLuX3/h5KHUzcRtKJ+7V5DHMy3PGy3tyCfp7V9VT+j3xEUJIo1hORcpOF
KDvKkvgR0SdbKajXigSTAVn+Xeg+G4HsJgooc7ProUG2Z2oXdiSX7fOq8AMCtsH4yEYUUSBkMfYQ
QgJ2G5WaYAuvj6U8w+l4XGK7snVksV6/Sz5YD0dK02+QxCfwrU49EMvQUro31Bc5ovamuHtNDnu5
e7/Qj5+a8RGTi2RwoZtJkfA4EFRUqrQe9KeqgUn09SSqqhIEpaoWjjrbqxFyQZfgN06//gN2862e
qRTPQyZcqI0QEeDCaj8bmXP9r5HLoNZwRs9wcejBIlCx6ye7jkqfLSN1VE/tge3RZ9txmspb6/S+
ZsCGCvwHUGu0K8wdG+pe66Q9VulhHVGx7DxkCjprq2melLZNsTp9ZWoXrx9SJxAhimaWcYeB70Iw
BAye7/JEE+I07T05RaGvKeKWsWXi3nA8NaBZ8BiNztr5I6BOuSwgyy/w78ThnElSVXACHGdRBmhZ
YfIXhExRVldhJWsNMSSulfn9Gw0VaWdw9DohYekwFG0P58Yzhp4hEEllK61dAVVVgTt3HphA7elO
/W0za8hq0XyvaWUFRTux3mDb/KdTBi4QnWc7CMNCr1CuC1J2S6JRF3k1Y558tQze5aLxu6f6uyDP
4eMRp8Eiac9+B1oyRsV4WdntYQsxzFGyx2ma4j8+O7+GVCqVtPmDcEouM+dcYN0sZn3hOaejrr7l
mfzQ1v0R7swJyxfxOJFGytaapvb2nHJ/zaEwTXUP9EP4GsNRvouEUcHozatAuBD10Vzuq0vsCVv0
lSJr8DUbl5FmvZRTRuvI3seB0wqRMxwwOnmqXbKYiPE7k9A0xWRUuMxeRMxwVoMDfeF+cRAfXS+b
j4vZlVbauYw82WE2uhH01afeq8I450v/QZeNnQl36dPffIh+xm/Py7zoE9SK+chZ15sx5KoFcb0q
tluqG7+OIvJEzPwpRWxM/7laVbCeACAEqt8effMLynMfxi+T/NRSrwZMR/wZ5aZq/UtU/+mI3IUR
XamojCpyO9qhS6LwUlE8KofShaR1FwMBTyL0mQDNILNJGzI63QXJrTZaYw9lq9VBvANip2cOLQm8
miWnTbDMR1gzTKsYoyS2ZBO/y5+GbLlfT1IwbjIN0HfBuwu80Xhyoss5sBDvwkkgH6m9PPNeRObG
SUpSz191aeTIX8jKc81EANlGTj5MsAmhJYU6skZGxqXlQi2P0+Wr5hzuct0uV/NlrGl6mG2D8s2y
6pEb/DE2PlLhhdDprfhsSPVzDGgO4ZN5szARckLbXR3PUA7M3MOlgqA+a7YIaUIeQ9hrYuSriJKW
mgSJGpcVrMJVqGmLq/f3tAj6lPXXKi4IS1tZfIwFSahtzXoA3yE+gVMzEelH2dmVIMcKrh1k3kjl
2khqPA1il5a6Qz7oWW/vgRyjysO8zboFZWEiuxwffLugBfLmjbgNuw6S8pP9mRUK050uO7Z8cKXC
MpO3wlXiX+h97+7Hb6FSEo+cNxy+RxQlr8MzMp7gxDig6FQ4esVFd8//zp5fc98BCOoZlSy1gNwR
79x2rob1Pe3WQXYf3FE8+nyD+uXjTsmUrKtYxWe0G1DnE9HqO+oWS+iTXhGf8tKKZ3ZvbGEjLbIx
t/V3HW18d1PlQMfMbojm0z5ViR1MSv5hEIPH5YmbjaUMaSaNlwuzA2Cp4XtOAhPUd84yA7p7xuI3
NZ/cWQJ8jgtbgB9iYY/mcwv+OMPGPbK2PkKKFv8TIZT1FRHJ6IglvMlyUY/Thfcf9E1PIa/XOA4j
H//AflybyjJdGfqNPGIRDPqNWtDrvcsQddzKq6FuEEY0qov3MIoRqyxIjytgtNOpNXmoYs+xOI+R
FjbOJw4CWa8yIW8v+7wqnvWLamXzEj+LLHJROQiG/zw/SiLYV6Id2OkC+5MPmibQhCFcSPEksqS8
6KvJM9HDG3rJogK0Np/qWm3nQSUng0dst98T9TJYCu7wnwGUWvTXKV7NZXwKpcXaZL2uHJEpbId1
CrES9eEOPBfoQ6CWwRy5RaUhW3LevKRgr5CwCBbJMSNxZcXEX/qrNeISZwDYa6UJIyXuHZazGBkS
DoMNkRTxBypEAOJ3klKwsTlri0cfPW5uaVPWtGL5Iqw1TYt5hzWJ0DoeC3QKBXmhhAoTebDx7J7o
ILt/0hNYE0EExQcccqVFEYAdG6pFyHGw5bEgE6vwpXZSVSRfgSn8pE+lEMo/5ejvNeySnlcRs0+i
FyYZgWmBohYtELhlGh32Ww2M888cLDkUFawl5L9wXVUaJBx/dsy2JbV9diJK6goKwRE6smdK0vvV
cCZnha9IynYx3fHJHNhUYdY+mC3dA5B7CK0Cr+eIt2j8BqaucrdXKZUq/5EufVea1up4zvW9l5Mx
TTvG9eGV5RROh0RRtWciUWMHjQttH3SfwM+m8Ma+lfTWEfjacWueA7Ag3ek6j58Ec0VIHJxBg3tF
RHmEwh4Qyq+J9o+obukCuv375/EHJWA4Gy7NW/x9CgliSAWjZO/u35LEx/iO2W7Vlk1nhzxTdSeE
l1RsfNgILILwumpccRaGCWljfFNgRIzO9LRSat5S2eymCBdpfxoAo3Y8P/BrRrTIaCwDhT24D+Qy
n8gDAOQPGTCB+qqZYcjVwJQTnubQhBFV1UsPqwsBV8dDtwpi5UjfO+9gR5Sr1ryZqLzrdioCSWAf
imVQjVrmXfjP+AvEL8tzMoW5uUcNsGg9H8XSy8YQsn0kpy+FZUs4x5BC8T35ppEPtWA50K8eUAKp
G3v6mk+YjxZ1HstsFT4iEiy0PCpND/TranQ+ah0y5dpsZHPyzkvpUfgUXGlMZvr88lpr83qVmBD2
TBwcJvJBAPgFf4BQoM6q2WeKAP3Xl1wJEcCJ8D4Vg+BFD2Z9sow2IC0uq3bqM7g7wdscI/TRwRLf
t0po/6aj9mFZ1NuNe6tLab7xe1raL3GBeVXa0aIoIfg+5bWl2cGtEYaNGrshSKdqf7zXuHtZh2rc
CPr48vzjuNJvjn9xig2YaZt+hwsAiBE/GJxMb4UwKufFgqADawp+UApHeyjoQZr/p3WpF+Fo37fO
57GHBIFVLhxZinEi2ISMB+yI26DL+uis8BVksPzSJe/jmoIclkCg40eA9hcQcS90wDsSFIuXrYvE
QbhtjmWshaHayvQtHTLPsXqwVj86zmnZVLXWsiqrGbQuxu4QC2JbmLwSSnMxJVZaJkgrNPhj2nV+
Knk4PM2uyFymyF57VVP+PnWl3rfQzHrfns2fIC3/DAhUiSqmSVBavgsHH+bxIkkfSdMl/NNmhbtg
acwmGW/JqOLua1rIt6U+/zFqxYL1BpIy7O9l66IoIiP1XzQmc49G6j2tKLGtivXIvfLlhi5eqbb0
nZuu0P4SpdIrbcCbaKCjuP0Xuvm2Vp9qZU8hL8/FO5qpYIBgkpkFbecwRUgs0LtNOq0vVUsw4XF8
BICW3fPcF1KaqHwrce1yo44pXT3vMte+zJ2XhWp5FTcQ2yXPOELM/lG9gYmWanV7LZ9kOYrqUG3v
opZ2FNCAx6k3KGGm0CtsjDP3UvOmw9+c9+8Jtjkw4wALNUnAuY5mNqeul2+Qvaa0RD1KSSKpka2V
YR8MRpzZTd/n5bKqoidyBtvwzcDUY9pwPHOa3XfTiRIWFZUd612eoUJnusq5r8hsJe0tgbRZlLtd
HDvm0CQHTinGxRWfIMb5sRVfBLs4Sni8QlSmJLem+67ctjQ+b+IP5SCib5D1ijnReQVnyz+/evKz
IF0XMhxC4UPyXkcDSOPsDpbS8B8j1B+tQPbrhe+lDWth9U/zytVaJVy6TkgskcHnEgBnkx5+UyXq
62tlWM5ezCKzpQxLJlrayocrrC5dJePkZeJNTmBLIZ4XX3NSciEraPc1Goj6BvUr7bDN5qNSi8Xb
caoa5UzWXL/NBbi+DZaYMmb2M7SFoRm6z2bLg/dGlKratlGpuv0jU5lAL2z5OgoUI2u4ycjLEZmN
goANqbyWqQj7XCL0gnWIgJ1yZcIvoKzxdh5CBCHfAb10QBP3mogjQ3UlDueHz5RtI3uPac7JxPoN
k+kUXcGPkJcXwsZg2QNtb9w/Oq51NSDNH4pDURrmy4UABv0MHiwaXrXnIqRoXPjZ6fzJS3dAhjBU
HDCxdhebZ9986uZc9eQrSm0Yoqns0KNSAaENrBDD8K4O/PZvOcyjG0cxIQL49dHXvjZzDvIv5f0m
1fb16sg7ecaZ1EUbS+k8F0LzqpC+4tIcBel4KB3CiqS2hR8pYJxmwSB9dXoW/LjKVxuemG3r2wjs
nCv3UMc1dlnjTW/UhqJsd9UutrquyOl+97MO2aiLRXT0WbnOzNasl+ar7ORyFotz7zCsAdAvhK1m
ozb2cC0w1qaDVpy6zpFYUvC52X9o8xNYs8LooTtftY3uWIEGC/GdwLgyXfqBJE8t4qz+d3rXxfYw
wRXIy7rvxXu0/sN7TnFJUWofTiYeauq0PI+zS4kMqNfxXodG/X4fvLqBoGj+UMMceXWtld9a6Sdx
w1enrguDCCPDpPZ3EV6rH/fu+qYz38wdTR1ODzc9NjnU4DmLd6xBJ3hdUZZGCmVUv8Bnqj5Ds43R
Vs7bFJ8wWMIjp9t53sXJag+en9hiGwHNAZwtdCoMbrIvVBoNp3oXRxXkFMuZ7RikO73fDP8Er6I5
FwOZVf7BdORs/58HbdpqL5WKja8Fll6zigTy/GSRbc02ijIYOekli4ejTcMdQTK8hMe6Kf8aVYEz
4sjyRHmXdOpC1huYPcH0p2YoRSKBfbSbHRriwY5e/xbzx/4H+HDwANlwQMByumhwz63iFsx5abP1
L5vJWhFE6mMNC21tlV5qA2m3VvqeuhyOXtP8isvT31e6+hekXBdGp1+UQ4OPIb8WLHgb36Quvuve
mc4M5txfXvBQ06V9hrKvMzbHMRwhJdL4EmHxk3c1j8Q1hLmbBQLC9aptHOKbGWRFsqqV1wHqPH2Y
iMvOzm/J0LZdNR4TCu2YF/oSNrMsLXAXsZFo8LzUi6of/1ev2NGeJ69dI5on1pd5MI0CkqJ4rQR8
tFLMqwXuQofZ3k+0KwnlYKnEiMF+96rql4XoB36sjvXegPga9zeAVLBonhzvVbrxtSd1LLIsvKQC
wPyjt1KZ2Mk+ABkcGXTuam7GN++Xqt1oY/HKdqkGR0Zs0Q1b0qQWV04AYySs06VB/gaC/K8FDkaA
9Z1PoFh2VPB2+0WjMxcmkyIoxQ7w9A3OINkOMiulZucXa7Nfb1IZ3yD4pSdDE3R/2j9Vbdlbpn6U
bcczQ9jRnj1gYIFQUVow7BCqTN6vsmPT6oBCzwHr3j6DEeBoNBxIp1dRzuqu6AeHlCcpi2dG+JSv
FKVJHF9EBgKB1DS+j9ZQaRk7Ssl5VchlpJnn+aBw2tjV+Q6BNsUhUgVZtk3G5DOIkd1FOb6zbgvE
IDYsmOn1cWgyE/9wszREfSSfWQCJ0WYhpdzwmRtTU1kaPAo1lCTuCvvAO+XGqYLzTit5ALNZik2v
qYBCAhNCXj7UJsgphOzwdkmqe2sWj1051PmOLg5mDNjPg+M2uNkK4c43qdyMuC7M3IvKNb+4QBU7
38k15qdOl6H3+S1uY1a+i3AxNuhGV1GXp9B5dijm5dj35SzZtFrYTO7xaCmTksdwBchyWKdzsh4l
gdQjMFahdy8KDUW9qD2sLj1jsFPiGlZ2SBRTmHH5z1FAOfhzENZmmTg4Vcc8DlyF3799LGXgrT+3
3TvPGgqMJh1CnSr05MXhX3Gd8Cn68zwjdfEUidD698duixvePvmRLfGPQxJtNxSQR7ThEsC7shm7
cTwDddUJ3LZzR/2ZZstgfGaO59nMk/cs8BNYQv07I0JRRk0yhIjiVuKwSd8/qJI9bn8geDIuVD/I
YaFW87LYSyJtem1h4tTr+6wZiGNvtIotteEQgh/cTsNnzdrTOKfL1KCWi9mUYHF4t+apc4f3mvmZ
rmobRXgAonvcZOz6uCu8zZC9vYJsqAJaIDNZzGFOnwuGu35Fx+dTn6PW24C/+paXTSJuMH0pOvvq
WBTV+VYdrM/MS/WOHhfSybC2EaDE89E+fqgL+RG9pyPGt2j8gtCQCSPLDNw5cURtwwqk6wCbn6hs
Mr3od/XvfRv0Y9ANuat5eBA3XkddxNcEkI3ouZIFkUhLZMrv/WGFGjdLLf/kiTjoTQaJS5KhR7D6
vt9uGGRrjyKm2lc1qo8FpdvpNhXipfqAfMBDvQQwY4bDu+ptToK6ES9vl+KOpVG2b3z2uWxkG6UR
vnZaBDAnO/LdWD7ytWYxsE4dJor6rTu97PzVH8wsPXtpO3zd7usypgMnmt5Uje52sIcmIovuZVb5
mznEA/7r/6JQv/RFlNEvmGErFC0YTrJ+jBUtDG3DNXAMDnbakqk9wx36UWVjBZ/NffmYDlqV5ARZ
iTzhgr+IYxAPS01iY04LFeJ6ZL/jlS3smIa6B2wVXCiUe7u0j7pn8pZO891rxNxv+0TPTRM7AkhI
V93Zb91PJTcTQZcfscPQNPLvIOcxWZ8eNzhs3OEYKdZPdSuhZtNtlPNmzhDvD6B/KPSm4l5jMw4z
zCj9o2AK2vd0RM9HhFT81JvpIOgAqUT26RDkez9WfGJNm5q0ixzy9zX248k9AcF79GezEq55Jxgr
dCCP/qq5sAieyhOC7SzZbD84gWNhWUs2AQQfobd2wlwRFDhbcfeDb1sbIgaXzBETON6QBrUIZx6N
gqG3wilSmx8mHOt5qCppRltNYk65BWNMVPCa2vdYlYyEue28mumivAJ2FRBBvpRV+1rslPjqN9b7
5qD+zOb3P50Ydgl0Fue4uf6Se19ZdW8Tq/aRb3jW8Fg/BrgAIHIGVfyzYSsJOcoLvpQCfgAccAfi
xE2qIuK1OUPUxmZ0W+5VluQQhaQfseeLuKcqtBm6h70HYwyeYl6UM54Rq3ChGqpWnItUgLIbUIuB
7IQN1ZhCFPoqOMZAuscNmEOCQT8ZxuEhd60ITmWBRorMhkO5Nt57o1i5BxLczF4wa7hKou6ZlAvC
8eL2Efj8DAQBqrG3jG64z6sc03DnaST/9InyqoXBnOkRtaZ1xl0w2gEvWC//tL7MC7F68hY2vLOA
EXk8VCXG3Whj+aQsVZ49/2ZuMuOoP+c8A+mcAF6mnuBEUeF35p5LjnEn6xvCK46/6V3y/1MlilgI
Lv4QBowr1eMDWbqaqP+XjToXXUQyB/qpczvg8Gp34E1T6EPLlD9xqt5A1x6OWyEKhqvkKM0p7Dcp
0CAL6K9/s1ukc+OwL8Ly5d5I2cmmMCjJ5WNtjro7KFPrYCrDuJBmkoQv5Q1mSrQaRPm97JRsZwJp
GRiqqHdXkjVTNf9xCt9JXXdQ1TsCHAX9I3kEvfJxJ/t04y5il9QizTosdOnQLKm8ZT0XDQEIQhJs
+lCqinxBxrXbHWNVimHZno9e27HSzDhkqjuO1TrOESrqHlfXfTQkIGywC+en2cz+N/WP6okpxN5w
pqpepc2Sxu3Lpw3eeZF3bf/6qeqw7fE9bwSMk4ZVLoxVIULspfmQl3yFLvks/PTkEbgloD0lNDeV
R3J444eT04LOTuE48WkvSO0QFdPsxg/kA3/Kygm7C/0qRWeJC97ip+F1H2MsAXuwkDPOm9dxDOb6
M7LBbkcvLaPQHvy7MbJVvljbuovmjGtxkVGmtLcrBl8LNmjORLcZ6wLgB+f3oE0jeN7XaQycdkBw
zuTxmCLPBEpriYSyXs1GTsfGfLSd7cORQRLCZLvq6GSyZU0A65KsydV4BOQRHlJ7YDDSbLUg9o5T
Rlyehfv95Wse5qTcwjDbvJbZhbJhRJhDf9iKZ2ILYc4trAsQ6u3gEmm55+SE5DJ4XStjIoXx7MSv
f1V5m3yQutgrub2HQI4cbsBAc/swME9ZgHqoOJK1pzZGrWXi6iIAAtXzERdAwHy+8O5v9QLdvq7y
1TGWp1j649uhiWU00IraGH5HFgmvcK2lC2BGCpfN79AVAMlNq8dkw7xcu6MdlmCrtZT1L+rwNwwZ
0rP55FzbpmTk0Iejbgdft3ZIlhsijNd2KAj74TnjpZx3TUeAbeCY91DcvSS1FT2TBdj+vqfmWs6Q
VjkpaYFp4JT9ZEqZ5gQrJjErhdqhqIgdh9kXrTYM4uwRZ4NCKWkcGnY82aglenaQ8epNDIMk+P10
sbtYcLBuhdBswJBwp70obKPNo6HeMw5dEi7ISEicOvwvPY4PD7Obyd2q+wEgasc2jLnOuQR1Fuwx
5UycyNbMnt2pCc9IpQeLr9vKkdwumFbPw4enG3QYroHJcAYO2KjIVcNbBvKr/hMZwnbFqM0hwxpT
SA2hWwRNOEKOWWt4eWuq5A+JMDt+TDllcWl50VgxfqnOAR6EWgnz0Vwn/qfS/Mx5q3ykoQWkbO/v
yAckGEcBQ0AEF+6zcQlt76CSJDCPoGEvsM3VWuyHTWnwe10+B6Hpoo6q77hcfXjgJGHpCSraXldF
ax7YxTPyxgpcCqsw4uT2N6kcPE0a/mysBxrQZIIgmanhPYkQeXUmar4hsH5YASUde1gRapDNhQga
9Q2VI7FZGETf31fO8J9F7NfO17fq0QzkHam5aGJ2VCPXCP++9i/7T5MGD+dduZvFfGEJIEKLOvD/
MN5hOGa3coqLnl1C9AkXHohlVjAnn0evsZeZ9e6g3T+c+VtylozrIVO9cgLoDeJuhzc8UpCbtPF4
yMFAPg2ybMbmiThr9HMYX+6AQwPcRk96mY4wYDQ7zQ+8N3drjtOEqfbLrCRZLbJOCl3yXLjpSJA7
hwMIE2FPqLdehdtsGS7tvxTA76HkWnJ7iCeyMzdf6pShz62pkSOfjTavO+Em23xQ9N7A1gj/RDt8
CeDESPzj5XaV/HqkGNdZEjI2s05xBlQyq7lt7J3lqtmw/Yj3RZnitsJSnVjFi3xALU6vCQrnPZWl
++l7oaliosnKlDa31mpzMCD67XaNK9oTchekk3GUO4NcdGen1otBiaWoyOOmJj5pcT0lDdWiTHWB
nh8rfLwvIGg1EEk9qeyi9g2xAjI2e8lJohV4UeSN8kOg6GokCfSL0tgDEgXgcwEfdEF9YULGt5/A
NujJ9l2Xe1jhqrMhJqcUcdbudMFmnROom8mXHuRmEIrdsz8OwmyxmLntP/AfG8ThHfnu6rlsgqsg
5KAXIf3jrOaueeE1ieiQ7h7udQ0cY5fiKHzshc8J+h0QHnDiaDfRlJqWgpL86cOW052z+4R1BnsE
ifRcZ845PZLjIb96GFWw3VQvEXtEHR/xMxAGGD+lSw8HJIfh1ZkdZaBpb50/DIa9cD0w7AZOeEia
0cstemoF9xgYzm6ultVqjFgIgFiAdk1SGtjvnAcaZcENAHn91addvr10jMDLTc7g2oyoybHQA9sL
qsAedDE2pnq6aP/P9qaJVPteZxtMoi/ymAv/usBGKDKO6EDKs9ep0YciJKdgPXhQTpK+Kg+RRx6B
ujKg11vqewN+Dsr3bFpSPV+AHp/hV1oqCWHUxTmdQY2TPDb6XRPHWalcu8KapkHYQa4Ds9b5m9Rm
xdDanOFncZ1S+wH5ad1qDW8ZdyhTxYo6tL2Ghsexz8/csmkPuZfi95XBd1I3OiS/khaYHeFHrKVL
gymQvqYGV4i9o9OH9V8+WiBUlyUjoxEumOrsnAyf/tKIfd11MWxAD+jmt1JzvyPOt0Gj7ah/VId8
etsCPxlSU7t9c3lDks8yENajv0xuF3fbyNjrREJsZV/+9XsM03mStVKnvDBrvULaZOOnVrcGrjIJ
D8czQuxPrEErOR0b/s61oH/crivludsREBtQEH42KkoaNLh4Pp6NqWLuTv7LcG57vb+6pJ+KxRSf
21fIwPCwQyB/uqx5Qf82WfR9UNdD8Gk+lqSlMlOQD26rjFerbIVsYWsCqEp2vtq1Zj0/RROcdMZ0
rU4C7r6gX9l9MSZ3216WfRFdAH7xZDLoh3hrA8vDrDGl8uur1sbUBrD0+dW67hPnY/i1q3Peuozv
sUa9LrC8OMAwWUvXQaOtR/xXetZoDppsS0m5XkLFwcRceYKWUIqE2ck9a+wRIZ+Zkhw/o4R+9loc
eI4RGQGprEQsWZ2ZCeueNzYhnwHZwXFIClbDsVV9aYFUiA69ccV4n4aysmgiGqXdVppnkO7MNrWQ
1nDcTjpQsLXHD6N7CpqVo+sUMkMGoTDWK6fuBgfeUCjWOJw27NyzZVruWupZ5Qz/3WXZ1oiiZ20G
NaREPQnC1sVWgUDhEJCyvzjwS9ON1VEM2YFk8UzENVIbjslveEjWNOoIs+N0l9lNtnPu9E3YDchb
OSOjdiQRbRkm7DCh7aoPNRegHou9Dtodj9me12hnv4eFMjUJ8Vla9JTGPM86UvmKusv5eibAHrTe
rLfrK1E6XTCjUPlO0uMMU+i4Cf14UyPXGgstQR4NbmTjOJK0KrpnnNF1s+Io0ms7ZQtQNlUU7zO0
zzDsT4U0i7UAljvd9iwg7gK2dFvb7FDQ3YpU9uuq/6PNjUgfvK8w/TpF3f7s2yjpvV6f/b9mi+lq
6B2vb6iGSvy8w5L/db8wPchEoy4+oeL/i5SkUaiexEqH1DzpNC7MeT2/Vgco0tjyAvakPn36QzGj
WcPYj2DxP3GU/NH3/cVMSvEZg+bEMe4iidc53ah8uVCpIWhRGKy/nLUZkOBy5IwW6F0u3hHk8nBg
W8O3TnkpEoDqhZoanLrCYqaFibQsE5dxfMZfYV50iYi8dTs+dmyD04UXDrCbgHv6g76py9kNu0TB
cEItbQMBwBg1956obwesOd4BGJUf0SyP5fJUxjNBxzUSpyL9B36cEU/osjRqdI65Q7G1QmHi/A/6
QflIoNp1pghOHdrEFPK0bo0ztGRESsQGRgz6wxsiS1Unw4F++82ropVozLVT7dg6HRgDwEgLU+at
EeG02sK/7CD3EDmmB7b6JSfhpBB5PjpN2rBCpFWheJ5jHEIdpTcaK7wsxHj2YK/nXzlsajgHebSi
EN/YqzHNkFWwXa5rbKocnIAhfeJMuiRf2PpKe3xSCwV48M0avemPHKB6lMAM/GJGx1VXIkeZR3V1
sf/srh2Sco+r9q9lGPKpCGF18PNvjbM0Sqv8XkeqU9AdQtRBXkMPLCXCsaZTFRl4FZW3DmPynveR
KBDHyf6b20LqpsOnrT4ZcmSgs/w298tXVomi6eFYCST8r1BaJGOitUmwEyTN//v6iAJcHbLt9CG+
Srx7RI2ijetcrw9pJGp91WRuIgSaDLgz/27kwO92pNJT2IrYzFgcKvg35BsP6SVe0opgLKWnzDy0
+1rEVsGBX2m+9ZYqMk0VNVxVkHlwduAI7xPsUXLu1IM/cPCykN122neZt3cNDOUCoGjfDW76LyAE
FPZGHR+rxHv6r8P1CY6j0MNnJtP4dWBdk+4H9t6wu5htbea5CmBjbB9e9oJk+d0e0A7ShO5/1seV
PWhrK5dZ0vgMdfOg94fNtrKBfMY3rPkhY/Em/JODLjcPZtvbYYMfw4x8uuzlaERP3Wq7fPWZp58f
jcbCMrH0sDLmcFcWNbi1fBUidSdLh/2RgX7xTuA/RsqqXmqNO5GhuhF7cyb0igBMj+gYXp5dGKG4
OhUFWFDhG7vKBK0KhjihmDjd05uShGxhMQhy88Rlukw8vpqBgopuo2QOT2JpY/zaddKlNV6rM287
cVpCXo4WvxNHN9jfxCDtwzyoAuzKPb06zOt3ahGUdBDqLZMVFnIbEeAqRZVksEqXN+LokqZcSJyw
JKZqd+C11+Mxip7+iPRpIJbtitbMa+3NufWz5HihAMrmoIsr5LqeiX5grSfK36nlKYRa6ob+BMno
maZmaONQ2tD5I8jwEZkzIjvZ3jNXBulgytFWbVmPLtNdnH2GsqKLkLQ1B0IkAUxoP8SdJe4GymRd
h/4Sp2M8giPPE4wE+Tu6Zn85YLVrkA1yv8o/CtfklkpGDT3AXpBpY5n25Lu045IM6h9ulPTU63uL
cvHqHcHTFSVwJ+kvmaWDkdPfp8jRleTxu0WTyEVxQ9Wz1jLnp6aty/Oy69/sAuvhLbo1ABBp5cza
DrTFzvHrNANZ4ReCGT2TqIEbS2950R4gxro4tlnB3BEfRkeZjbupGxErCIClkZ+KYgixdiTwX2WA
Ok1bDPdxcEhLxajm6PdM4yIe0DgT0XAZt4i+pf0+tdO6k3SGuUwInv9xfNmdsuYaGZg6LuH0PB+b
BFPU9dDzuhoocRCBPSn9C3i1FNXc2J6nwjl7Zll2OFdVRrYsil1bMu2Z/W8m3abc1CWqsrzEGQzO
1OAmeYDeSaVjwQDYwblWK0yFkuVehvgmm+De4ziS4AQwTAId4faNYaIAQ0G98staGf4BrV4bNoSE
Wus0wHvHW4spAkx5KAypkbsOef5dApgvw8R51tVC943CO6o6tgfxV4sEwTcPKzeyiDMoe7kB74xB
o5xtQF3yx06Hp7NxAN/rEmYJUxTwMYYfMdwINktA269LRlMzWS+bPgO4hBraFHXFKRjig9+r6LyO
hTg5Vhw9wV/T5J2vUjWVXsIUJHrZe7n2Wt28djVW4ksx9y0mXjktrfqOiL5jBgPuWtcuUo6k4+Gw
CbGtYlLyxYTnSeO4aNGv9mZ7QthcoPCv4NiE6sdvThG1hWF6uGJ40mOx7CSXBLh/dWImJQl7V8fY
jL/iY6UelkriysZSuL+KVPzQfypPT14lKbvB7MLwstyEsNLBMHmZoQ9tyCzP/6n23keQolvjNsK1
T0AoEHc59VNfD/M/bkeoLGQ4xTs4N/4k6x9niVyfio4RhS+urppw5ynVOylwpd49m0ldo78lPyL+
8JZa6QWymjyH2k2BywsFSnET6LpC5sJeCam4xdxdl4Un88GJwWojtrD6jWqkOjl72iMTl+QkAryX
h/c50DoEIAkECFdwNJcpSsMXVEc9+ISy49qE8VpGlkF3ZGksW4K8/TShk1/sKdcIKp0+PYDvsPVV
2qlCyIfJ4jOnh4vRpmrU9JxcZnvknH/VWqaHsvNrmoNEG+A/iCDIkiQ3I2AovUkc5dMSxjNPQRR5
cqWe8kBox/OdlzEsKZwxzw+2Z8Zs+xCEengNha4ShX+f5omdZWyn9g/NpNcx9mYDHk3cb8xH79sB
MRLRXbnZmfsBvMbLWNdkQFtPRwomrNiM7k8cuOMWo9swoosTZ+nFg1rPcYFXCnHqZY5SbzRX5cjd
o0aSoVeLY4Jm1tO5QYU70maYXVpuvCZrfVXMytAmR5wYrPE+cHq2Qk+MGudDvlc7JitG0aFAJnd1
hsnZbCJi13CfdlOGGipAeISs0NuAki7K717M5U3SYswR++gQJPEh2U1Ks0vf5xGCm0bfJy8HMbWp
WUCpE/1XrWXbZjMIS2xYVQoIfzCwNuX1JFyER+UXTRzptiEVAd8gqNYfwHhpzI2zRcZCfd3Di0+G
RlfQoL2/D/Uy1/JWBbhoZcYKLXNdbFXoXXqaVxnzRi2fwP0ixGpD2nCGx9vPqyBwJ67ZglBZ16FQ
5DVHNUBSl6wn4hcAI6psi1dLr728fxYK2ScGeZXgyC2900G8FPj6rQTSb6dx125O2CbPegxJL1UX
yZBYL6c8GnBM/tXWsbV8JF4lHgH3aI/jPOQJ8+zEBmcchVTmjmjafDotIfsF9NfPZ6y56E8xQyq6
+H2w8FhE9T9dB6uzsfuNrX41pzVSa5voqmMMBEf9Wkm4j2MoCWl20kF+u5Cx5Qswfhjn/S1EVepq
rj2ydet5a/aA8NY1wNO5pFwkX6hRbTRmiqSWGrVH2OXsR/cFbc03pJp35WaGqBm4DUynEyQGQym6
CaTo27p8XNSH+iLG57lClWrqWzyhzUdrHF/JQT+qBh4bUbWrZ7lxUVx0D57MKjotzL1svuE105CP
gqKv7kRvQ2yQPG7kvFDGtWUkdzN1DSlgnbRuTQTnVcDP3vZFpvcZoEvbOqfKapPdKgJe3gTJk4a6
0DhLnE5kOxzAIajTfJzdLvgJLnBUNSxDMdQiqzjd+1XezzGRElzLqkUqhqPWBGr+AuwWyMyIx5hg
MXDCjH4b5PaGDkwY68ne5CkivGSJEJDFvFOCIrWVlOTXnHvZxV9eN2+T6Vy8tWAKrwto3MqV0pow
s4aUE72lNDgxFIn8NwUEy48Y5c63gPxCTVHqr1g5CRrwfJaA9OX3OWd1ulgvqiBuQkR4Wrmd0Kx7
lKxizyEc2MwavDpAjzzM1eHjMVo/KMCE7nCdjob6xKSchrS2S2gY4z5uzPrESw4I3K5yLM/vUmVn
0UAmBKYsGr6Y7RpYdljOf/wPzFQhf8kWX+QORvYvaE0JeNnehEEG2EbDB4GFLHBW8MecL9pUUH7J
dSbT20VfvajJif/4yi/uQ6d0FrP/TgvWCNxBQK7lVir2upmDdO1vPuKU9w6BB9UOyRTNRi+whB4L
4zHlz42wTtayZc9RoCUX1EOuKCEDSvV717SpjgRudFgbCneTZhvCLVTalqOJd2qHuWeZpl9bWJPv
E1WLHBOi93Dad41KHgKEAwun0CZzbwP1JO34DIiCorJmjvuXwh4ba4tKD8nVDJ0kQnydv4HfJcul
loFC1lhysRoTzM3z3XKvaht4vWg4ZjfI6S7iINKSbEuPzype2CDTr33rhvBwQU1N+c5gWBXftTLl
6Uvx5Erf2QmXKeSeh4ZX4ZpR/Wphq7sjP/Rmc1U10AjGWfwyQrDYDzZutw6R/EAM8iPMTRQe1XTM
XxSSvhc1GGWWkU+Xdow7r5NV/zT3n5eknyusbE4/sl28toSS7P7rbM7OEeGwoXVnnRuZbi3TsapS
EHNFMUu+Jcjmb4O7dymOTE322IwF0YnQpej+09Jm1ZK2wLLmD7YnPJ41M18Q4N3rObLn15/TcJEF
tjkaf8u1o3sq+kjz5xpfRH2NEZiQQx+hy4kLoeKoQSM6xJIMWSV2jJDAP8+BxRZuHeBbnqw2Upz7
J4wj5YPqCb+QP+zeBq8SXEA2h9CGLBlX53BIORHJY02IiHUBuMfDjwP9oMNTdmFxfPhPGl8S1Kgl
VsVt5tFNlSYi+x/5POLSvCGoJXONB1w+RPLkMuK9fSBEVTMu4AWv4TKioTdY1DbAuT3d1FcbCk+/
eY3L1dljJAH3aIVxt+1br2bsAwzAWQdDfHvUeqoSl1myp4sFC3peNdknmCf+3wZHCNxWict7FWcj
759fI1sE3mEwqPW9Rg5sp60QHdaHYm1epYTHPdRQAkoVh6bRTE3DjopAm71c68NmD/9Z4iqX/ddL
zC43G5lNAE3uiHxnu6CP7eQa4AUTAjDLLmCnS1kDQohesGq6JMnkbPo5szOUFtf/X7luSnw2KSH0
+fVTB0Yj+YnKG69MmduzO2CYBY+BDym5li+ZneKLTybTqDLJs1rhLZ3ez1kXNHiPIhApmrrXtN9+
FQp8x9R6QJeMr4rIszm0RQhFagWXvSmdgOn2fmSHm5eLwHBYT06XI4iFALo7Fuu09uXTC/7lejAH
hYdLZXjef77w0eZC35gIzJszvHl4F6SPgoEOKkgXmIQShrRj58hUqeLw+EgVKiZkV3Ik4NnCb+oq
NTvvj/9sLAMEr5lwulAqI2x9uohNRBgXyFYDG1+1PD/TgwtvNSvrrr4vz5hl5GpeCdYCcJiyXJVo
OZ/w+kC//RGmf8a2Tqvh/i/XOjpWdbc1RRvFkRNp/O/pv4CQhYFm3NrpJcYBBKZaKMeL1Lwz8fKj
5MT/H75/b0eHJDsegRWckLLwD0wQry1SjX7BaXD/whYyP93gtnskXhcyMrcgFHGz+jugUx0Hc/Cx
pKlYodXc3TwJgKwwUtt/+u5saLbzRlpSLkde4o0PhT9ZolSntEOXy3+16xzJetdt5q3gJ9fl0wCv
FmcF52Jp8O+GbKo+1rVNYaj06ZtaKR1VCKAXdFeXbZa2+upjT0eEeLr9CgKtKSlDb43LbyBc6nmG
rUEC+Yw4qNCAenc48vn+mmio/tQhGLJHhsqIBVTEUuIS+ckSnzvUQ/GqJ9PbfGDATc8VKmnE7xm3
tm9vYtGOov3NsFm3kVqKZa5dYt33MgiecZHFJFyJzB8DfaID4DBbJbCUsd2Og0tMruTmOXW+2mwt
e1ExR1dQ+Se4rWw+XiP4g7vc8NW7utF4dZmL+gMWxT0C1ZpB4HCUcw/UyFBd3FJwjcIfMywwA+yZ
PXl/qOZruKC0NkB2dTpngs45sEz9OoUDUMyKsj5UCrLcCoqDGzuGiYi1eQVYUBLhQCOanAhMf0Vr
vbTAjOV5yxYbdggmxhb6OI2xCxpwePswl7CiOKdAlRZCHNnB4g1OG1kcje5MCLcj03Bln1Hug9kq
FvUKqBsWIZ5rwzoc51Et2gI+EdS/HuS4xE1eMfHO2rJwM8X6L22ly13kxlmum+LljOiKZ+nk1/us
ICyq6g3RriAjxZW+zVzTAd7y06PjjB/ANBACUbeoUs75W5hmohGZi3XM1BvBuGM91RUTV2ua6ljJ
14V0bGYmA2lkdjixl1DGd2uNWHKkp/DDHZDHkb1gwh8oxUuhI6K9R0gV9xL70tPWiSlgIlGVzoB+
TmTTiNUaheUQUHdkRBKvRYax7YnVooV0foYw+xP/aWHQdTmtRo3sxzogutknsGB+kHT+qZnKNg5B
nyuMlXwYnJcShhwhGJfhkLNg6A7RHA1oXm/AoDrdXSK/rrQOiE4PVK2+sOG+HLBuksJmsdp/ix4n
7iX2jTAPBv6Os6nkNR6VhOvT6/Ll7oh1a+jUw12LOkewf6zjXv/MJIEtkDktPseSPoixT3oaXWhm
Mb70f/NDEFXJb9hkvkx1z041ocwTttSolTSGPeXv/nwxhW90djT702i4Uq0BCV9otG9XoMvHVEct
RXUye5mCmoB3YHzh6KA/KjdFfIUrvFBCVZzebqsvbmhgFvcyXMkCH5te2P1/vQInN2YvOxHuLAA2
OqNSr/T6IiaY0vp235/WVY3ObwVKcyYvKoc3qUJqBUfPD7BUuds45hRVD42hG1AdsQv/xjF7Of7n
MkSKnDF0ErVspBJi6ykHcXmDRInbL6Glr09XwSNrzljhVisr3YOZVFQNc+BHUQM4da+fysLsAfki
5A3AQircIQdkC9SKa7+kvyNXc7qKZiATvUPcec9fRStYx4X6q7dpLOEDnkndFYm5axJVku+mYqPO
KQgdFDIbT/LMM8CDWm/HxvReN4bWhjiMVd0yaN5nVpGdbjO7YIcDAY2KRX6/cZlMZbHAZ9dWRw4/
yPwJh/rajnGupWWfhkyYize/meLUl0BuEdTG4nIbMpSEjFSkA+/eKXZRM4tM6BIPh5HnKylL2UkB
dOi2ya6FjFOwaggN44xSxiWzgZYNAGbQX0R0wH9y2F/EIEh/Askl7h6wY6PvOWN4EmDl3NrmvrwN
jV0eUzB/3NoG2ojj/WTBjjyPmUlhWt0eNwnp8wUdij+tG4BCdZdErXl0HN+YMvgkEafZ5i7RAmti
PprfFxf26fM5AD+mKIYUrvlcJSjcAQ5ywZugkwwGVeFgWaCNq3LWpRTJGeXLFpnRHXP3N80mD9wQ
b+vdoP1zD0GCb7MwcXJNG/uEj6M2ubODgC5OiW6T67YiY3bdQ2NRx3TydGRQOf7exEBM+Wvx4la1
SFyeKKRWOJIot7+5ncC7w+C9bVhjqbNNwMpKCgTGZnunLG97koCjowKYsDBdN8jvgNH40Jem5aZp
wwkgEtaYESZGvMWWyARU5EJqFWFMtkIIwBLKuaKuz/hEMv5JhbqfF5fCXimJKItJpfbcYmiGEl8c
3A4RRz2J1GpNg3AvcXEmvq8AuPzEMp4xb+j/oIR0SSWEfFI0p1nVcmIPIGValWGkYdBl5L/RFLd+
S+ie2sf9rxPU2hGk4q4MQpmFzuCnYnYki0NE9xwrksKgpvMO74aSGw1pO9za0sXQp4XsAdLV0xP4
R+4C6UK2DMcKEWU/W3cR1V/DSOnelhRfv2CCFKiZkdwclJMwIR3FhZsBvC7JqujElaKDDe3ytsyo
0IXV2WhO6yxEKGDB802/oq5HNO/N8UzPvKl8QjY+6kE+0jWTtWtj29D1ZSwiA3Zhz2SkYKzuEcqO
jiaw1//m1IalXlpiZd55BGDomz2npwXMgN5UiVkxRV8Q7R7KD53Ck8Dtve5j6bvtt/Ks+cAiZZqT
TmTg77JarRo5pM/GBA0nPgFpinfuwmcIepWvwH/gPVzIn4/gBFIUDeTMNYDV67pUfzXzp+8+TDaU
mXN7UMTTuGPXPJtBkq4LgPh39dp5/UWBjHcmE5oQCCbb1+l183usNpGwqpDG1zU951zYdYFRLDOw
klv1tpE46rKqg+HQLHh4G28EkalD0dYwuIXFVRQM4SM1pM+YFf5Fh8IzA3zz1q8RJ685RKI7JjKg
uYZsypoO6B5pggP1sKZv9AHuNoWj+RReREvOa3+a2wBqyW7QftG7kVf8FuEYuG+U1ecOKamoSM5O
sPGZWkJrPpW42bpb6Y7S3Zvu700Q4Ex8ZzGfqWLBKicRA8uKlhfxEGF0AslqyfvWs2H8bcujm8ip
gz2y0YLd38K8qeavvWyIRvBGn34TkKqaC62NW3Qy8W0AeiLvp0pNFuUDrc02qh7WUt4HIENKG8Pg
GyO+KqXnXdGPbefLqGhOgfyZLwN0BnaCKWtwvxRatMzVJ+lVmRMsm5LSh5IDQUPfCLzSW5oTTBL3
OovlvzP1LK2zFiCxgWpuXITsX8UyOP5SXWOn3aS52cpeMk0rz/5n0pg51Mf09zy4x+/eswSqK3PR
hpT6bBkeHQbacdfwDUwBxHTG9wWEccgCbjsKVqeuilRv1cH2IhKwbquojwDu/c/8aHmQxKugvWxh
SGcAzNcO4wGIMyaPqHLskkR8qN1l3bE4KsMd04Jw1g43zC0ww/TijkYY3yz1DUxO/mNKMjPItQ2I
DtWX0oMA+lk+BSieeyX6gMK3zgAEtq+CoalvZrqppdRMfo/khdETmVZEhiFVSKS7r64mIgrchlUm
LmzA7YtZAkLsdqIxqqkkLIakJEVm+FHRYpueXg8tPFbGJ9ZBhTJIm7Rux5egrMAJeTRkV7WpPP/W
Xrb9B5LxuL9mfphvzAg9H9aVPyDeH3mbVH9sUPeaVZqQwReTZ9t79IMO5x77XTzAfdFN06eMk/Wo
gpkT0KJWG4v7DoSEiJC/cF9ZHz1FKPi8dclt0Lj/81IW4C5HrOyBp3DQTSg7F54msMkTY1x7ir7m
Od3Txw8ZpbzxxwyB1MFg9UToRYlg7wei9fl6tMAtlUyWRNv1Sc3dTP41ElDuFGD/3Kic2dcUIVlN
M1+Gnv2F19aSSLCCyt/5dkIIW7KiocjZkxfHkurWDzaPWM/DMYk3K0X8cTQCPqKYQnEjQVuEG7Lb
4q+oqQMX3Ent5OXlKUjRwTZmjNyc1G43NE1MzTjZ878qCk4JluSMr81Ala7/DKZ+yqQkLuYiSc4G
GYC1WGb6xbUzYxnCVbcn2+IGTrXK9iXIz8/v6WHqv/mNSwbnOqEjBDMBebjTHlnUGW51+HITay+X
Qeg6VIQlqdfOeoQCw9hR21fBXbUVmI6lZbhOh/hT1NUc09+0bkd6EGCqf4KYmMMA6CS302Ih8Els
1F6jxcQ4v257Yzcgkn1jQx871pZw4YCZO2B/wukfA/f8m/kIPtz9NGMaBjX8+0Fj0R3bEtVLoloF
T2aD57RixjkttOW6ECvvMT94fbJuOo9ZTAj7E6zgVYhzfrVvJlBdw/NAkFmk4omoEwGmIj142v+m
sH8a1dwbibJLWf15kjyO82+dRs4TFe/4BX2kucGBDM2/+cTmkf2gFvfn+SA0cRX3t2Qpe/HfxwuJ
gPvFGTjngBGfiEmPPEl2QmwthGiUAcfjxWGPMCmA45hXnulxgjKjxLMdj01iEiQArPu7K2gcFlDy
GLiy6BYzteqLMbiuiZBfF1Ho/FgWCYeyeHlbeUOF3pSn+K6pXcuAPlTW09pZaMa1+EeWKovgnRsl
avclVgNOvtp47QtOxdkymcHIHkxZO+ZV7p/Ynmam7UybyDG4Owp5T2SCjJIexI/2fXzt0O4FjIQt
2GN4YQkcH0pZDbzinbLUMXTe47fSW+gKMdyjT2tDFemGhl1/M8l1qlrg2AHlG4W9XLLzP9xpGw1F
Z8VdCyr/9Z3TioNSSplSSqsh5r08Kd8/sQOZDG5sFGe9QVW3oix20g1CoHtghw2YDp4tSY313GRJ
XnGWOmJNuupPUwN0ttXt/V3X3pD829uljqbjaTcR6loOAazW/hyLY+HYYsyXbuslFwEnuPV4fmvx
rIwIH8g9XHblI457XUQjCJpfqiG8P9Zr2d4uARPXKsZohAkiC1gezUDTK9JQ1edilTH151Z6hrzA
rlFF2L6YNt18V/13NW9Nev8MpwkoFIEIRBFwpOxJOY0CZgRSR4Of/4j5a+LscsWhUUgFt0XggNz2
srqkvNp2pdM3mEY8xy5vWwrB0v/1FSBbfuB/e73I+LkhoUYQ7zdf+9PkkDZ+53gTGbpuuvf7HMEm
geqQuH1bsLAyoD+b/mhEnTIcwBHCx1YYXivZm6j3ucI4Fqdhqicquf8rtaKIjfX/vkOqX4062IIb
JYXCjc4Txc7PtNAP2VwMJwk0bnRv6sL0gKsE1cRiyxEIYP2raTgJgfAGZkcncTWvRy30bpQ/uafe
z38uoB5aOovQyoZcKmC9U+GvB7GtdDWHhsgMVk8f0fxx9dCEw2OvhR8RH2F5hAHW+yFzbkgZCwBr
UTlaJ9TbLWVzVNWm1+CHTCqRs6oZ3YZ7LlizC7U8keeo3AGK6UhhwFo/OkIqCx16mcsRYsvdgL/l
VvmE2gUUoPjv3PtIz3zW06/vCRKEMcmT9lfJJMt0CEzfoTRGYOCSZ/NihHRHKRHFfrndQx74wYfa
a2O7ZH3LOiANiYfus1YJ9jf3zLTs/TktYDpu+5rg6EG0pW45xVX5qnzzEmCnPrKcmonjTMJcbUty
UiOh1Bj1QH+8RyfDN1Dtf0F+lN6BDR/LPjA5KOAC8ay9sFlt4DO+Q/acI5692hQ15WmXN4hz1iAv
oiI7uoW/3ald8KRLYGL+okjy0womdkt3xDJCaKDXAfproV92U73nmiHUA2gx48Ukml2SqaQGaeNe
nLFJ5U3oaz1s/95KiDH7TG1mYgQX52S29oqZH/ieN2pM3tdT4o4vAREm6T3z5ESZaFYDOPSR3vhm
R2e8l8iEV1ITXKZ4uDoFR+0yQz9R86gpCDfsLqghLCFSLsm7PCqBlNerhrYnGf9EiUa2rpKBuTrp
m01fUfTunEYgPd/ElvCcQ9qKb5a6wqRcjfp3IA3bnR7C5vwac6kO4pou2Ow87WBQtBqGTnvpcnzx
q1N1tuCH0InmzfcAvXG7AKVJrGPlmn+nUvH8njt/UTT+k4+0S4tX1jatDV2UuOABmE6ARKB1yCnl
YtCqOI+gyAHRXqFAn4XicsC1IvoOjMkICY7v3gmufWRHcYq1dHiFfWkBiDKnnkyrOdkhxKkP2AZr
fGnHMQudzsJ+3H2UiOer5ZoP5QQoKHLULOm6MmoY//I4D06oV3vTkFupm2rnL1Ibs0R0OrVNFgnv
I+L0Fy3tdXoyMPJf90JRt9mlyoT/JjbfCinR2CxSeAxRgBRvuPoow7seoj6ZAvWhJ95axzQVfYyY
Ue9hz4qD6hsuvKSxSu23TCnWNBqwUpMf7hnjvVOZNH8KtLNAJTj4wagZbK4buqfnAEf/k+uNw0c+
/tDdOF53bWtXeYtQQwmiKk2wrguckJaKPndZeD7NChdum+xFgm7Fld54OFKAihiUW1FdONlxAWUx
RpK/EfQbIrfwORkPglwfiM9WH6u7HHkqC5Ozjpi+o/HjLSpRsyDh1VhE1ibNd7cN9gJBK2oOIDUm
SrQ+GKG0CVfdZSnTYP3zNhm62YgwxCBSOkt19g6DOrewCHnf+N7oBrojbtQC2iNi5xE+nswUhgAJ
PYzFDs1sSxq4EErPnosV4vBe1hXdVDjXofPdZ2WZwD2g/b2EEMoeZ2cTGMK7OWg8wpOVNWEm4wRx
qWrXUr62mV9Tq3MPbCoE7o/ALbd8DAt7l3phTIH4gn6mkZbXLO8qfka+FNYUXeflluFx74kPU6En
vAojubSYcauEFsr8lxX5iCegUynTr67LC3NkDs4b84cLSRg9gC4nQ9L7f7mCMf1bMfdiryqXMtz0
3U4M8ruBJGO1jc99zX9T887rqngyFjj355EG2kiZQEP3AXQNRd0oVNltgMl8BW4rDmd59qs7THuu
gnNudAuqopTLb19M4X/wV1twYi6YM+dWKH6klm8YBZUTf4bJpcHEm1OOsJxH8o5etkszM5Syy0Mc
VQGxcDYRfFTEBNIiZAmRTokKnQQErNNBF0LBaJB1YKrj1/WD3qwn6T80UCEhgJc5qtO72YFj3XCK
kZS1SrmxehRozT8nl35WUSJ22X+8AN9c98JSmUB9RpmC7eGubZac6O3YIbgRU0sD9wfKnCd4rcQh
B3OZqH8+EmrH0RnCY1pZC0yZSpqYgREoNKeD8cXW/7R9AsPkvIugSr/EiX2Io0HJm3Btg+4k2Ped
YCK3cfzI59+47FWlJi2GYXLWdkwckgdx58x5u8F21Vj8mUu27KNrQobSS/zXKrdzKQqxsH91/408
2PwBKG5JlxeruUKuH537LafEb/zuENpztHw8OQi0izujtXo2H/OfCJf9Ls/PuxrwgQVwUHJ4UAKW
CHY+eoNyi/zXZ4WQmWa7rluypL+7WrvaZfl4928Y/DCQpWzH7KWqPR6lXk/JfxAeBTkCPkYYfHRb
jNh3yC5t48UnpIqQv1L5Mj2xq2cUDtUenTL/hgtGPFCPF2DAG7eV2KpE61kaHIORhwMkux1E+Rua
zm7kpVVV2yIhA5tbCgRo73mSI1aFCVlWNxLci1JD0TRYCDl5cKfv9USmvfG4YN+sS/DSBfyyjswe
3M51zKX2MrTF4O25+B2TJSLbEf511TZKz5tw90v519C7T2BFMhdEVos20amBj8Bu3i1hj140nCCO
PfTYNFXjY0Z9wXgxa/gfdYOCidJS8Fo7GHv5CCk78VpDP90o0H3JKVvb0IuemAwdJX5MEpiCHjHa
vdYj3Thii7anCauCFEnso636EhCjZvvdr99YRUZ3uFV3bRLfGKs1iOkEbQFXcAcmkMQsGbdNKFNP
LBtdsKkWZBif8IrSL163EY7v67oVS3uD+Cuuz61V+bTA/gg2sK0GBsRmh+cn7cI5Fc/NNvoT1edW
Ha98r787VtoNkjj3CMrUH3yQdQU6rm9GoRCavzxKOrEzV3z+/HERE0ErjcQhfItMYYnDGOd3suUR
4epiAfB8DA3Y0iM+gzF/suoW3dYyR7ZjoXgK+jvgSf2zovNIRQEHGCYBXUKPlH/cLVpkjRhmHR7Q
DuIZqKs3CgVImeSb3aANCyZKE6dtLJZxUke9GvWsBwEVYLiPsAHJNg0eNARPvVyxwVrZZ0S4bvl2
xb/y1zaXvffStEaPTGbn+iwZicJuSiL+4ImTXZnqgFER5v2Epn3sUd0O8u+H0+i6aOgdbvL3M8Lk
B5WIKJhwZXPZjNZcDhtZmdPnNMoe8mKHO3Ek0CGz6AO7jd5sb0Usjnbzy9qzND/Y6f4piKRbW6U9
7y7UeTauFuvFB4TrpAHucuq/wC5jRiytEMxXRNlsk3vKei56H9UuZPXWZMEQ+2Ac7PnNG8CqaZ1l
sJOhnsmK7aQV6jeVLCQWAbgrI6rWiJCGhVMgvm2TavD0p/YddxfHUyNE4I9ceBGY4GXW3R0bwbPC
psB4Ihm/Tfd+Db1U5I8W+uRiorGhRAf+lTdeRNqak6I86lwwRTHtrhhiwu29p2nz27Q3IVemTPwU
csMwkPJoCqwm+nZ5Iv+erRdfEniNxxl98NqBNB4h9VKv4nGIOZuuOFIvCko77r6BXcCIsj/2XPnj
jZTJmkUD7iB/MEiEDuFYe+mZOLOTaO4+UgEBVGCUWYV//ABALcDdBWlH9phrlF5g8yZmn1w4K0Nl
mO7ApLvWEKayTU7vIdGQU3GsawD8+5q4NRkwFV3mHGEKhll0O0SmsfxnistAgL9L15Y3fGMOSPdB
eRJwtF+YWaZpkJolJzg2GFpmTokBegUTzPHuQyUEn5FM9Z7pVcVWD027XZPlUmb6g6JfMAzRWLhp
MBgJNuDmpLDcTxg3UCb2YUnU6vZZXHKhYhZEDkfB2WVXqV66/Xv6wcR8yWHFIdOibC28GWX62Ipp
yf4hnnw4cOT5mGvsHfYOTSgarx4WAjuniNDr4sgROEUn6t1wJfUczjomhDcuhn2+H1YA/JkGWNmq
d1ZJG5U6c/naGYlGDMTZiJXx6UAJdp6tMHlaHrhb2aGq4jwwhAfRlYPffisnek4pJekBjGPHm2Yx
AmQ/ENaVX/1mgMVooHsK8V3/6cmXgb7AxUrifHVXH52oeAOQe51/qXkh23iChNKWRT8yxEv+tmgC
b38Ff0RT+t6zrT5myRFC1hRjTHi3MbwtHq9YageTkS4ietF0zmh4w2QJKMeBxa6FJHdZTfO8isQQ
y5ZVqG7jD309pdYFUgSZcgRfkVX/pv5NgeUho1+EmMd/3ZDO6F8z/kcHF+nG72ZKwlCY8Y45TfKp
ijTqrtfZkt99RmtpuI0A0CuPYRBTQriVFF6mGjpCQGPKhje+y7Joef+NloiBt8mFlyAb4FTa+r5t
HCBoDYH2/EHYQEYRlq9VyjtCdM4LJ2D3HvXr3NT6OQr/gUFrPjq/0LAXnDouMJo726BX7vxrJXJC
UZq6SZ2RygPJsM7QS4YpCkuH3OlY3VrXf+gdn4aJ2+5YqWGD17nqEWwlA6fRKlzxQWtjxZdXg2FP
J0WM/ZSsas5dgcayxkWNx6jpbqy4GKjZZkPMjDvCNbv4bF7ePID5684mvlAZgmuOJ/A0gsXdXQqO
D6wHnYMRrTgf4ospbaaORVrEYtNY718Sqq1+RY1Qu6k/5qxl67PWk1fcIt2zrYcPMzar1Ek7t5Qg
S4xn3L7mnt04X1umj89FqQyoGDB9pzF4IkSZDXN9TNDqgI7IB2M+jh/HD1NHoue4aj6BvLRVaLWx
h8oKJL+LQMx8yrgZXSSHGRPLCQwaitgkEc7U0HJ0CPz5wkXtr+a3qqWAtKi1iuO7NgNV8cHEvhKi
XAJqcr3xMe1WMesmX67woTvLephRuXPZjTTyDBVt7NIdoNNoZ/PPAkUT3ZgsNaiSeU/WXHDHfVwM
zNgAmGXl2GDOGZvZYJhhn+opCghVJu6KrgXkmYrifjRGowmF1o2c2NavSqdyS+x+tfQiwfV2p12H
GMl2/+iJuLLb0JoJ9+Ariqjs4INmOWSGUw2eEcAEJztuo+rlLmaHFbYRAUT9f3VW16j7duH9ZPQf
jFFPVGfITdJWRzWtS9UnNEiqoRhbN2UiwM7/XoclnyUxyaLeI+JoDz1DY++REaCuLLA/EmgzpFYV
dSN3SGdI34XfIikEdgSUTy7sGv0VKGxEDT9pSgr8A3eyKGPigItEJP77vu5gCOy1hUzifPfSUm1f
UCNqPUtYIn9z/x2rwHQV8OAfehzt4zOUJHxRsZJicx5bk0WEw4nXy41KbGwgP339ycvI9Wjw4cib
l6aPnJ8v1mwq+gLTnLDtMfWPFBHfrnHPqPXt/CpCR6A9ODmuBmWRbUocg/p0FZVeisPVlG6qjeDh
fHBQdHtto6PY53ABIe69achCoft7hlR7VqD5EufvtZdFOViclMn655QTRpNeb7Gdkzg1/Hp8dvU9
Jxvfn7MbY1nMGBF9ai8aw1CNxdElymoN1wSO+XzLYvJCKeXMeLkHCE8VOhasRWOwyAUwNOw28Pch
p87BoD2j/YqWP0AHCOUiAcN0Bv2vi2WBTAJIBeT7vTeXPXF4LsMsQJp/vOeysxR0+EANXtRTQWiD
DgrOzEVbotPreTQhyocT1El4CtDXA/jPp5dujtcWF2PHnW6uZdHBGGvv53bDD4LdUHkGcU5rc/Om
qnVy3sYWSgXmgkZUdtqJmzohWS7RraD6Q9ZiBH4Uig7FgG/R+CbPwKZ0xMyCRdg4luYOoQDVn4Pr
aHUybaFkTeY+bQWXp/1FE96rPxbRqDbiYygC6NqE2kkQTtwx4+yP1lrltJzzp0XQDBGvW++A1o38
QXAWEBcuzDwMOwQj3YhD4Iy3u9DvqFrx9RbqVWPeH3y4Z7u6JrpD2399MOzUzX1YoDx1c6yJOwyK
yS7yYCBALXzotjkgm8CBHVRgelWuQX14F5yRbM6wmpwqy1ln+r/XepO7auifdc6XsDI4REjs4p1V
eJMh54m8YgaY4Nq7VDlFVZJOrGHwiYv2bWv0TObcspQnh1CKPdujFRF1RTL151rME8F1YuisqjbT
Df857ybY5K9dx961YMu4YDjUPoTk+2M8ptR2R0NG24Oc+SXkbdOygiCmuxLnKvWCQ8xhYGydXhMH
ZCW44u6498L9YUsftB7AWdVjBMIne/GB9sRO/NSp7/6raedrytcBFSOk87wmn7py8/QOPE9yp/D0
CxzWfA0sPDQzn/tuaYGWqW+lHuiPqtHm/yS/60lLAtVRxfJtKRHpeWNY3S6cQyAzonFwxQGkhVPu
rseAC9WIEchfYJ4mrgPhiHhlAcV8H3LXLYgMQCJpie88SQZfPcDDNhROb+aw73kluzukM24hdkJi
zz20yUhu257EEg85EfSnugtuP8OwesD3bDM5dvFVVGqPhQJ4TgfHtKAoPh6SKsB5BfuyTq/SFSu8
dBvUelRYW9GPIbZeIhsHn/60oSRPkXWoKwgbMnCvoP/GjlUObvrjhQLtPu8qc/moDD5ycYxrRxfa
d01hjXRDVPMtlGLT7ELedtFJiMH/FcsupWjpgucwEwlaQd/8nTj/cXeDj+RsA5OthWkyEo0IiopR
kQl3Izp1108xJVoLZ7UcuCHfWrtUCcDPrbBNsUMEbAmRbW2DtTcZcfJUHNsfU9fV9P/cBrIQMpUG
HhiGy3Dg7MW9mJOlgEUFyq36wU8YkhwPx+sogbJd66MSP3//DGuHWEWBtP64838ifSK0n7n8jvwi
nTsrnxefsREiCUXEuETkfsBuUP5CSWO334I+UG/HNvEpEa2FvqmbGqEX6J5lqxCobFmBJMZtxept
LTw7jpmd0ReeHvaTk+FQKLJZQ7d9qMk9P8qQV633tsqNdSSVIQz3wjldIL85+DfKG2jaV3VBcPnm
Q1YNe5J5u0sFDpWwt/UDOnCO92W/usgOkxw3aLhWeMeVkywj/lLP+Yt1TN4hZsWQmFkX0LDsyAG0
503a+5m7zz8PE9gxCsf/vMgYi6NdrV4FCKIFskp+p2Y+VRWUFMmrNeymvyGaQuKJO8nmDYvsvIrj
PlQfnAfEkoSV7nqP7QV7qZLjUlIswF9wSBfLLrAOBpu6u8lorhNAJ7tINgJDaKLVLQ83f7sEV4QW
lg9DFjEed8TsUiyAcNzEb0JgOm2iIyNv6gkrzzzS3OP5dWTAxNEWCxCYP4CTN351KWPN46cjoQZZ
1CCq9EZiJlzznYZpi1+Y1ikmgTxLdZjOKwoMq3U0YMnlEM+no/xEyhYN1EdEN+NXB5nJmef5jCY5
141icw1ZRxIfttTkeVRql4DsoZtMWs8/QhPlRpE+oI2LffJiAZ6KUOXC9oSKFk5o90uLL/Bs7x8M
qOvyjZiBqvMW7SglC2/h92q73ABl+7w9cuYFLn/rnJZjoTI3/C5shQY7lrtX43WU0Qj4bJ3D1qBU
9pgjvrwS6vXTWgHzvsjNSJWwZZc6n3j6muND3tMjbcjak9IamD2U4Nr9HzNy5wed6bG5IHg3tEXz
SLGzjSGpZLXOqNhhbQggDKPLhCTO+1cUriaGk1eSpHCNUVGBqe2WgaOJ/evL60BhMfsKQ0pARIuW
diaYNIsMO6gSYw5LpwD+Xz8RN97Nu9Ru+cDwwKQUmfI1RZC5Hl7Dga5e4pcNHv0kv3x4pRjp2mSO
EiLqdAAvZFvKGbTxJhBtn/C7IPVSd0yRgqUYocU5DpOw6Xaj3g3Fp507QU7FzttCvRz4Pc/Wyy6E
e0+EE3TkooLhMjQqNKKKxD+a3uSwo/BH80k7W+o9B8GnlHuBkLkyqeqty3ZUUC8xmsNCT1Y2W/VN
7hkJsLuykX+GlJGe+MT6cWdsItlZRHrEt+f3caR/CxlnXdhR0NsmkZOGd0GKvjeeg3BSU/KrMmsy
/nYVv92LsICwiVM8rAvch4qJzHmhzrpNlyWHNfX2iSKNPSuvylwZhZ5ghxTzJ8ReD7X+afjYbNg3
6Xi3Y52e9e/pvEIdy3yw8yavhEtTB/1IWkMGqQULDdkXulAssua6VUtD9hzKp1RaTC3a/C4hQpqN
VtZmMDuLuU+yCGgJU5AFLnXbyzh4M4vrjAN57ozru1Pe5Z+X7SQQGw27jOz3Cxe8MtlFG5+NZ1zX
4F2tqJw5gNEu+42xFswcpz+nz9JCiKR+vXEUaR4/OfvKLH80Ua3auVTytamTIzkNFX/9N+NA82eU
zMHFFeZkejlcgK5lLsCSvNaoL0bnxwMihIjy8uaz9xIdU8N/O9N5iMjlsKVoSvFTZMzKn8t2kOFf
m1GOJZh5GvN5AyQ23Fi5FklpBSVzeWkkL4QePKMyoosf5eIAeNsn7JtWXovjtuH2iQek5um6pkUs
rJekrsGygNtRyBnY4uwWz5G9K2FeG1cW3pcN4bOzC1qvOvBRoS2CHL3oJE4JjGjNV38W/FNlgyeB
MjWkI2cc0LdjCBcg5sZNrRR6JjjqvpqPeY+Fv8QDa8W/XOqZgwKE37VvAVnnT7B3vbaLh6lh12Vf
f+HA+nctxMt7aTivguHabK5M2WGKHmSo8VRlH1sbiS7+emxXRFXTkYjXeGoAVBg7mS9V1lNlOOs7
jBAgs9nyMBuyrLLkxVj4vnamo++cPgqy/TCO12SNVGjfE31dD8B9oYmPXlLQP7kBvmjd9AZ5oVCI
ptFISYHjfAG4zYoZM7ASo2oUWMJdHpz8GlS+NNZd2D7bJNTTFZ/RyJANiAqzjouVgIDHVqjeDq60
TNmgIn8ra0MeM0czIXe7lH8yg7prl47bkKnNai3LYDS/bQ1PhGZ++uOi0QUCyhkKRDsElGpIjq5F
x+X0hxCwJ2EBUf8AkTtNWKVz2JLYHD+8NvNO58WUQVEzZwRKcm6rNCbTq6a7/DmYO9QLVCMWsiM7
bv1WNZ4jU3m55YFNexQoXK1s3vlaf8mAyJhzQGkAxdOJs5XKcaT9SLy/2qtxxMAkrQoTBvrWX07j
4w18kK2YOsDbWRwJQzDm2h+qOzjNLvI0+QQKGYuN1XwXJvRDwANiPOQCFnOzv9MQeP8h0aOBtaXY
kNWofG8h5Vx6kC9jbPAtcR+4jTjwKssU8nEYs1ZMrU08952fMBzOKNu5WfTB0vv9eqK2BtVLSxhW
SYD8JvrwkaAJZga0TLn3XJ/ppQmE9gyPETN6USnuP1uICNDUpbWPHhHFHIAsZ7GHfRe8ejaKvkAP
V/S/769rQAz8e9rW0fzJpwC5hn7OK6XjEOGVCZdTM6H3aahg+ccHdo3kW/HdCODNXFmgfzmBRi6h
tyh04xIguggG4byh7L0f3VhYFKN7lzL0qNq3NRnU2x0PfFOGRCwQHSLuX9F+FxYwPiZaGRWRntDG
DFwg5w6WT6ey/aTifgbzgdNKkeHjBjTJieSB1hKhH8/X576MVdw/ZDnGkqLlGzuE5msKoeJw0T9G
eskYQXRghcy20YBTjk7UnPPsihho/PwU3DE1+JEL5NtfxhTy+5YSzthm4vAeP7JfEIhbLvEAj9cM
fK9WwEq9rgZ20Xt7KCzQJ6KnBwlU8UdMTiAEtupWY2b18YFPLVPENVlKZRcJ+XJXqMHQgSZ1GSSo
B0wcykFvMtW8lnKos3soLzek8iIb0d1B+AUoiDcQYADTGNW7JzBSwTRKpSPa/ufYRpecqO3fxaxv
PFIBtdakEnRGaE6mW1Oe7y3OfpNLTLodkaielYtZ32tp/uqMbCNOg/pTu3pHnKLIUtiE/7vzQw20
+XjzSmSU7XRDrSKfTNhn6rYmz6BGHHQsu4BFPUreLL6CynVbQJhZjymMqAzP/zaccywmnP7aZhQs
ZGEyyu+Cz1eNFWlGlMWa1mxOLRnmwMY+eVu857LBUkR7RAPYQZ5S56ooBMeuL7VTDc1mj/4ahXpq
SxsReailY1UcDrrfF8J7wjgGYGexG6Q7Ux+ugQNiFk19gPTzvVSFZHkZF1QVgwq2Gd3n/cBR7z8j
z3QCPiCmRGHZQCwppiqJ90pbrbmk/F3EV09SSGQYngsBAzIixqJKG4uXIiixf6hQvvcuEnLCWyho
zKeXkz94/scBESLFpRRihEqvtOneNbEnc6ZhGCll5jbV1xIR1SlDVARiQuvgHncMVf9QvNB3PaWr
gNg+Msnhl969ufB0o74Fi8iFpLC7iAA6L8/6wagpZu8nrwj9x2ptpagrwb17xQJb1Trje7/rUxqw
GlaMUFWvv0JA45MEE8eo+5ahY0fnrkHcW6GvRloDz+x1J/O1evFnTNjt7dXMnRlrnxDJvTyl+im7
ZqSUsCAfU/dV8QN0MbnUWSg5XMHZYlB/aAAEsePFqa9NMssVo7oMTnSWyf50jZaKEUYEHnfFBILh
g1fAq2tuWrEPeDhfieWT8CcywQc9OWnWMek4GeO6CNMRZGPdvakHoPHm1jGOIf0EN9gp2pPYlPVQ
twpMHRQC5Zh+KkUzP8bvVsjIKy4tB7ffLn3R2WzhyNvyku9tUBOXE45MSTZQJzH0IGOD+rRce8Cy
WTf7EGF1GMqC8vg34LWnB3iU3VLvNkIZasph+HN+h8Bc+i1/Imi5EBNxUNyzO8HjzrqT91mImamE
EltRRIjuL/7Q9NsUAZKgNbCQBbQu5CyMUxr5NCkb7sewtW9NIse/Nj3O6aHybDiowLluQ3t08G1r
su2Hdvks8Gj49JxELuVc2uqgVuPB00lGoUsarusIg30b1e+VOoZf4EDFVCCGaMpSLnU4Nx6U5Xe4
u4OeESB/nSuqvUKFRpE4et/wlUH9dTK8XB4duyXIDy9K+UqccwpE0j4RcboXZJ1SvjF1HmcwrMGM
e1YRm+WzOoOtPurgkM/377gv1AveiLaPsUKwjoiMd4GF6w9ytYocVOdrEgWMEuwy/Z06n1pHv2SC
Gl1/DiqfOGA13IxtG47v6ypdzC+R8IJQneifSGuCwykpe8J6v84F6ZhWeHAx8YKZUva+b8c+I7gB
TMBtVWmvVd7xvpIImPv9IwV5FjAdMJ4W3h93K4coCsCIV4kPI+QZ4mHVIFWPTJqFKOZonI9i415R
BJBPWcvXWgnUqy01Qc383i/ERJHReJ5114jq9xCdp0l8yoyoKc1ck6aCK7Uv5bd3lGRtoWV7RMa0
llD08DNSxH4TFNbmD6WpJZpoUkfVMQN2TGtBqbi8/HBq/MkhH0AGQYaSiAI2uZPhqSU9kEz9C3a6
gmx0BgCtCPHqzuPfBNYtOybT5nOk+5e7/G2AfFwMIpcmHMGZL/5S5ww+uEQe8bq9ZTAzSP9US5EO
+sfByDKFfGEbqZvN1UmNj/S671oiYo9KAaahwcBW0bhc4s9sO5JGmUwK9ibq7l7/ctA2vhSQ+pCs
InTmPBNrSrUjF+i2C0BKrYNv1Wx6FhVKrp7JJtzNyF4AfUE7tb7X4r7cW61azqXeTQeCJnbh4cMX
r3Pwh4eT50B83oPJCOsNDtuvV3oQ+40o64Yn210OkaHE8b2WsjSThWvDTxOSSykFzOgD55oZEQ0O
CucBE5cG5LpPkrXPKl6wnJtZ9MCo21CfDBQY9y0mdD8mUd+9nbrdhxIf3rikud2t8vX+beRLwML8
XX7SOwRdWWbDhmvxuf3rq7OHI8C9q9LnvA7cpuEyZRqdtZcnlr+XbZXGUQuRsVpvV82v6i+a8S1F
BX8KXhjiV+QASGjH0jDlk5DzTbecwAdinWFmrBKrmFOeoBDHfMw5QpEshufRif0zKIlNGUM+pLsV
3iVDMkYW0vomNEcUgV0+WZxYhPj7813gP91Dk3uninsWM4TG0AIayHSduG888VxzZRKRCR3T/Q72
DTpNEmw5i43bnBK0rRXWD1StAEiAa5h+Iosg64hI4TxEeqnvjGZA9yOLvJgmhsb1jbDlyKXsIaRQ
dKfCuofmtuTvUNFsrcFV34mMfYUIlVOcZzb6jAPliSmUsWhp51+dEpkyjT3vzhEXDueMso3+Grlz
BJ2XAFquZUhf+Q2p8OtVD2FCAt2Wq6/OD7B5Ziin1306AJW4Zw3ukBeya1JlQ95RUjL+MU0tc7rR
/jyT7Bsqn4TXRA0gXGRQFVSwzl8HCAnR5SsQjjAD/2xYYjr4JnksqRXepe+64uwp/6u5GzvSjniN
JN5Tc3ZB4zed+gggfYVs9UtoVezrWzm907rhJLJ/lvFM+YzCsofdSbCpem2C15YR+jd0YeYy6ZYN
GzhfvvKtnJ+mIV1cAbtqyVv2vxVeSi3kWmFCIyB0QwyqxgEUgPwm5Yq7xHFLYqyXnwC+0FfjZN2/
eCMo6/ckW937Eau3rb+Yj71jQIzr/En2xh5yvVxvBEVqyAKeSP1FJNDOBrlcQaKt0IVGy0znwkME
D7MgKnrJvDK+HJ0h0keQWxn3xceN4EruynKJEgruPEWl+dWlV+uMR2Fmm7MxDj+fb+myDtcnUoWb
Ye7uxqO9cc4zStAmww5bX+lOQuqn9xW2jY156sJ7K07Z+0zygqTLIdanGWzZmTA1nExxfLQz/htA
N8OwuSQ5gdh8szVGCsutxBgDT5MQI+SeU0eJFAz4yXgpeCMLCW1qeEf0ioNF5CkKa45GCPzzmm+q
lzzqYTDrbJVitKFBUSbChgTm9mrYSPcIgb1Bcws9T+uCgyjiCuV1BqJ+nZ/lb+zFyipkg9PJufXE
sF/qcWiVv/bQRPKqrQSQSSSGhWJ8hqGYApUrbqRiTpyrd1U9M62qANQz6nlmXF+Qt6tGjc3OLiU5
9J+eLue4GYam2jiMsHch0C+z3nBYDVvSb2eqEWPvMG8QAfJKYCdNMyX/7b+Kpt3BuVCHDOHt17Wq
xgYKhrfjdf1Qcx9HhG77OeCEsf4rdxwrDEn0AA8iwtd+Opv4RscfR+tujG/t8EBQDkYO6U/ZFhHD
HUiILYmMYkgMFMu2c0mgAWRM5AA4D6BSz3hDehAJyGkV6g+Yy3DeTdKRLDbxP68cOhoag2IMVY0Q
k6AEmj16MeuNkXTVVko4uEBbz/GyJzsb7ubhcuuBsW0LOVvYOYnK/vsFQCQ+QODMqtPdjc0qgqxX
lhJHoaSftpnILgg/Kon7IjHWwd/5G85La9kHY/Wxrv/i03behlO+U2I3XWGop3djHwvV1dfV9Xv7
2uyMz9k8JDTCHGRIXIa9LIePNDTIZ6TGGKrOFUdXDiEq+mPVFLnAgVzH+Zl2ZsV4lmeMnLZSCRjX
dZsjUFDlTYERiayqhZ2mNUzLMLTaFHfYh0M3xjr0tIY8AOKjuLalgepojEPYXTfo1PcbS7VH4mHe
v4nDmeiZFfrzrufKiW0JV1oGqWdJqAXStEPJwxSjHNubocw1Zc3zb2DgWcXSFmI1y1xpfMJqhSw/
XZSVLiRkpiFdmhEIObrHKr2zsk1nl7i49qCBJZR/R+9yIpOuzzJonmFqY0cGqDok41dHddQHQULm
PlpYEREs8KtAfLGyFJeIuhzW/nARd5dQYouFJEm6OwwyIEBqiyxJ5QiT0/CERNu6I4U/4W23lmjy
g6OViLmU69za3l9VACHiDxDia6bvm4SQseW2TdkrIXa89pUBFzDQDARs0NSudOzdyhVlIzUJ/atd
HwJb+tqAEEz24MabhdUdFY2BSYi0YpajVgPru57NcM5QgCfQJDlDvIAnWVSxrYKl2LiWOsrRvtIc
MZfyx8Cao+91RjSzAymFVsk668W/YCV88Lpdljj2c+3fFo8aUuHuYW2mHAGeRA/O+0H9prD1YCUU
fNqI6c0uTTBlsbM8TsIGzAJNKb9VJOVqN5KvUC7IRMgbJebZ5AGh/mycwcEo23SYDmSzMi8wD6ws
drk4Z+FswSp8Fko1udErelfmxHwrhKEo4G6eDKM9A4l7IZDEiK4UYrn51Wl4Fe7urAK37+WRlNGR
AWpXL1HESdDudhUS2FUcHLl/4Frb7+kfX/EF36BtSbLXtWovJDpral6HgbdfR+VrvD7TbbCDcDBe
eHhGlP5OEIgJoGV+76qhwod4aXytul0gWZrOBRMQjcQ5rrOC/k1jMLo3CHewksm7hnHyOouQYmkw
XxQK4u8kDHPbTJXbCnPBD6EEOtIQ3leUYnzBjBAWSjX06TjUKdgq+WyClsOuNChN9Kvag57mRuo/
EvpqJu18qS6iJU2bfMWtUxzd+73qmTGGS5oZcAQJ7DauJHSIren1l714c6XWOlrp6Wz45RWu7tAx
kon7UGXRgEH0CJ+3Cxzb76HARjGD/yUemUNszdCVCbZbrTNergynjH5sUwJteq3LVELh7vGainW2
NgcUKxk2JEUdTIBtglpPQA9sKGRf3YBJiUV8SbUAH1o6hnRkj+MOJK0ttA53XsQX/YwofFXDRwXJ
7aHWZ3KAwqqeqZg2O0G1srMRS2pnvHhfMaL2aCbO6d8fd+2039mXgtQaes/lMkSM3iFT25bFNw/1
n+oCpj/4rxtxIYhjYJO7z2vwfNWmSrRdqAPUXpVgduWUZHezKNdoWKoX4T50Q9Qh4dpuuSX75d0v
1Ypzq3trWtQM3jh7jrNQ/KtYbY2Fgdsm1SvzRLAhkK49SMGMRHysVQVEGja709nbpKDUqZynZBav
3ug7v2Aihuzhe9PLP4O8ndhDmv9wPJOVDD6Jt1BdI83YPWKZjTEdMh3dolbchAujfirNvFif6q24
iySDi7ABc/LGxa1PzHxbcyTpHw1oajHbbwtaanh0JVK2zRePzs5gurDkmFmIRZZ/AbDffGLXNRH6
DTbNxgrJNBO8jjTvJxcib5AiI0K8aDugQVP9ihTyNPRowuZJgYscNy+4rnqgnafOShSK4d5DsBX1
WnMgHhnGj7hmIdigv8UR3PBZGGsa+MZOH9e5skMdOT2lshIjVfa1vbrjfvmkaDC1cYy3EOJyBqwB
Tzs4CCCFK1SgefbUM+9TZ2GU/sXjHOFA/usNKCdywuSHnzHc0dPHMSr5I276Xs+vMwVKWU4DOPSM
meWhjAYtywPtBnU0/tuKct3dyWNLskwycg13HqoWRQOUycPd4tvNpV/Jw6hqKf641zDXnwCR0ZgY
7XjTlNDSY4lWnn1jYH4NiqgRbNc2IVcxHxkbHfPO/36t1kOhwxYV9ksWhivRu54NMYfTQtDt9/ae
eiwhsY0vqzHUB/GNV1LMPBbeHDLm3WzTf5saPH3xZJW3r257a+zFGCI7d+T5Q01U/7mfIruf0Ds8
VaaGl4FUbeHljrq3Z6v5ZADmCUqt9J8xOvvNXoMeBJrCubl3a/lt3GQ/dFUDSExMDeEvx8dsfX9m
9lgAxX0s0xzlLAPwArn0/vVI3rGKBG2hOveOFmelPUXFyFHGlF83L746o76VbAFXKB+2DTACwYJn
IZ303pDSTtGzyeARR4L8uvNlgj7mONwagS4EWNZkS2wBnFVLtgRiVtdj+bodbRU9WxrqjMYM2Ptv
bGcvkn15Sq93zloo46irJrnv2Ey2qFNzWg097FyJR9qNhVfdtFu6eP0euxkL3b+ZOA4FSIkaM7Nl
IpE5ZDYHyWCNkxcH3cjs0icAf7ziL2KGwWWEP1SeN86GaYSUkRLg15NIDiXspGjG5o3DCvMyzBXK
J/9weI+eLQBhhcGqrKlFU+e8GWyPWzwYyfyrxxUma70dVLCoX24g7efdtvmciQlFdh+YE6LX4aWi
pSwVAJZb0uVjYkriH7Iggd4pMyDL81Etb+LGYndTAYKgXgJvaxtqa9bfUmYELCaQGnJIPWmiKycn
/V8yM3oTIMO4oAZZXKV+txWOdhEJ6L8fBGdV6hZ4NZEfKyizPpI9mLzS8gzTGc1s4pLzTOByDmvo
wgjEGNyZrFzyO5MgP0i8nxyEvix9j0O7nZOjeZw0Z4GjayVStnOotxnLtKy04o8Siv4fnzzu+Wzr
OT/ZP0cEIDp/RYAd0TLwmLABy2CfqBvAuU0PdQJQxTS5qRE2MjdKgM8GU7HFERHIB4UHts2RVLhd
BaqOf7Bba7TB47YyZVF1+ThhCKRrfZlK4PigDZUpZyM0T3mquk9K9IXD6r/BKH62AIBF/5vq5Dgn
VK6Dn3Ej1i918PuAajMOuia79VWmkbuBql5pGOnU+Fi+qsCm7dqAu5koD1Hzh1U5JiF451foGJpD
YgPKgih0ed/CYmOut87kAYhdl3gVEDiuE6w/jxB3RyRBgk8XZWbOcBwWYtIdpNkucFw5oSSBF9XD
rdR0FeBrMFjcU1JQl33IzIqXrmN5xbk0VASGDFgzcyaUHAP8cxE3RJ6lqgs3tp9x1/X1rsNSve1G
XRmC0a1dGdl5eFPrKP0CvPzemBf/QCZOBiV0lEgNcBqAuDz7dAzgdow1xTwud00Cv2cS77xdLbZ5
IuNTaQZsHie3M1OrYosrkg/2CbjTpn1f7RafswD5F6BII7fZTiwQ0952PK9S/egvZbXHx/8//TnT
YpGra3FTVJbcvXsmErYZ66lU75RpfwMr+0Oej8vmRqZFZKvLAXrv1IKQNWbWCBRgqr95kJSlOJwC
mAQ5D0qHNUWSq58EFS/Sy0a4BUW+R5bqR6hpSIyIu05Rq0gTSRjzkp+/uTooaHrST+LZZQJYtIJT
4ucEqCS7n0eqZlAGsxEdYVuFs1jjHIlwZlxKdiegAYCp8dy1aLS1cp7ygA4fk5r6uUp3ebwZiRzn
exTM7TjP5UDvTadOoqb9L1MdmeHmM2D3YWPT719pK463S5eGe1GhSa+FdEPectWY2LxigZxMWemM
s6jmHMX7J3He3SpsIRimCCih6xOOaMeiYmmSpV1Ij5SacDQmj+LqdAgd4Zzdk2kqq2tGZAwvc7lR
DbuNLRV/uoO5nTRfgVVS6MLpCkQ81yoiJbRneWMtS6FqnfOrdo4/ddV2KS3TwL3thZuwqwXL/Sn4
YXym45mozrV8HqXoDCLGFKufEjjXzQSGyp/MBIXqQfh3raZmGK/jXKf5akl8wOzKXJFBnOmMkYdx
ja/lkOhHBKxgozytkKk7d8PbjDpSHe6PgiTAJH3oUr08BigKju5L+17Om6NB49tfpHOcXjzlsQQb
zuV2s5qbhjO9oRc7t92vOH/m6zGvjvQO/VoG9kMKTFitQu2ajDgXRDDOHtyfpXRURItaWrUybANE
NI0Ip+6M/3nL7odWjebnWtItu7dtBsef492rVVDpxNbdOZ/70lL9YVLhuEHVUyBaxf3HJlaFPl/M
IVA3P2P6K2fZn/7bdoZsOwcs8/Ieqi8dYQeqT8HtUPSQInBEWmxAA2hzatv8Yf6wrLs//6PVqUW9
nXTxbHp6B/kqv6msq+988MvIIblcpweAiWnG9AFMTwijlGiqHNLmw+ebIFu0SuauLUACYF149wLl
fGC9dmU8C3mc/pqzH+ufD5ZyggRSvHv068aeumcvLQr28Mrbo9HIPQqxG/R00ic3t3D0yoUgw7u9
bV91BzLaOGcOODAWg7vvzGHsB6QSxIUCKvsEYPoHQwOaFr7NcWPEgTUDQbCSkyiAfgH8MQ7/MYzj
+wvaLi/AsC6oY2KDxGZD0oBJv8jju5pqqMpJdeLdfP+/BAwavnM+YB9K89M4TlMg2Q6mrWKX+Nb8
yrF4Hs260kR/4zimFCiW4KOq0cHvHFjCL3Zq6IoPWRdjaGm6l267/SbibydspntdCT8kdzDUN9MG
Mz14sXm2ymm+CE3VR+dxG8P75nwXoyrNHJznwT42QrD50+ThpBQdiPWgzZSZtfB9NHFh2zzf1hFt
AQ9qpMIgen+Zek6nqkEshE7l47ERhHQZKDAcewXVABGxrn+Qm74yCckO2sTodNvZ2G0lM+bCcJXf
H1cb8S8yQ4QGvgNi9hPjR3Ui8e+6YgO6lcU9eGM+/p7OxSv8qUTT2lJejiMpzCZZrbZ84op21cLt
m92kH2uYAGLc1JCJKQYl3XPhOI4XlkHvK8gu6l0DanbZLJKmw9gI6PQuE0d62qDuZDw0e9J5LkRn
Q+JqkZdXk+Sz0qSvdyg1lMrScOTaDFzThZLnbfjCb5P7bw8IQvWFBbSWXg2vnJkleFwIdtaL8yYl
6FUfaAiH13WkjaO/LLnS34r98Rvh88YQ+A8Zji3adU9/eJC9q63422//UJliYD6HBFmZeWlqesQq
dxmVmQft2QGVgY9RM25EBapU6GzY2pycPiMx9p+8nR5lCJxRdno6ifZkY23lzYzyB5WzNIDaEeWP
bV+DtgzTAAzkXMxu6Eghhc6tO5Li9Q+XOwn32YViD2S4NOUmpBK7s90V30GtTH8JESMtOxHPLWxt
OSM0d8wxEsiwkomn5zYeRX2ayy0B1Y7ammA61BuC6Z5XrV2sIDcWPirWo4yqF9vUp1VUVyQVnX/5
Hjcx909gtgS9scFblZIs5DrqWokmYR15nmDChYP56Z1afj2WL8BHKbnTcnulLgf+togHTKtmj/KL
AB8oZmB/SPSHZc/2wlB4zNrB0escU0mIDaiN8dybSSLlk64kMpVCrxIkA1LVklQIC34+4IEotSqV
oNyQA+h2jlk69F0O5AGjs7gW2v/22kS7Zz0M78bUkloHzp41cJyC1Caym7d/cFtu39RBMcFqtlvx
psS3nGZbcB2IiohMm6ziLHVLmlVmxbbBpEeVpkp+K+x4rsNeCS7/latR8LzgfylwXs/Of3FGlpTn
D43FMQV2bBIiae6vfevHyW8jxA16tZSsQXpQ/UmRY/EodftRSaIXU3FPvA7pzd1p5Yso2H6H4gAr
d6k3Ml/s7ZwAgSKGd0UMQImEGxYZun6w3i6sFNyF9kRoumMh4c2bc6CJzyE8kgPj/xaimNg1gKJ3
qQXja12hcKUyyUKlEbttLxEWciyjJuhcv7gtfsvEN1D5bcsaYEgmeYk1EE9lnTSfLjCJ1kE9n7gy
P0qt8/5YMM0ercPceOjFDS5ymPtc77dxqJgnt0NLFzt9RDTAMOj4A0Dc2MwTcmvXQg+dI9Yoc9NW
4GwUWnD5a99f4FDp2UNvIhOqt+/AEZa58lCDSWnIDHF06RIqlvr2pQaFxrPHakJ/jMjaF6AEgH+K
Zr9CvdaC/84jEIIWKl7iTbANM9PRwt4ksYZA0PyPQ7yfRbHgmuYnlVYLL1XrRCmPU+a9GBocGLu1
VShTeDL1r2hNzq20KAWlY7HsMH+9Sc2Vq8uKL13HmyW3dzRoW9Se741srdvBkGBY+1GGk8Z9aEjL
ApFHNu5zccy/z8DqnslkphoHKl+dNr9ZLvjtDjIxhCs0CIy0Us9n5J5/Ld6CqR79hGItxueqvi+7
45Ycx9z+kzLYDx9Dus0ZA/LTt1udBH4QnCR8T4QDEuZ39hK9aLWWv+oYNkZFrERlVQkdhhqSVTjW
/EvwsaEiuSzenjOvR930F3OxPwOrlLbY/IvO3sBLwU9O9bE8qt280qd+6IiNL6jkHCwyGBEqM/18
+Se+qcDbmUw0vM1PXelLqxrty8hUkO9/++i0lebRe9i+iPeIqDF6bRC/Q5txJV9vAg297+nu/lL9
uE3FPlo742RRNJjHCYdKAgQ38AasRPq7Hh2i+CFU4gH69KbTzHFP8kNIxKZivTyGdMN/Q02XCaqL
FyL5gDGUnix68+WfBgIbEic0t6NU7W8/MvNs6bIhp3LBbzEUg5JwlTKNKi17awQ2Xoi14YeemLj8
KGmJnvNF3trXkQNkrfaC71Ed+hTHndFk0ojZ+ASrNQJmyvA4d8TiJruv3TtvTLTfqeuPmqEVSNXE
t7tiCJJhH5BiFMldeGCngIcbUXbxB+nidJCg3dT1oTZ6mJQg86GeE8/+8LeFG6HzTpk0w0JF6xMH
DJtreaDttegAcBf+YXPWV+XbaYgeeZ6vIzt5Nr+KHkiMLYE9TgAAuDxbFLfl+gekCc9ycBGK6RGv
nNyDXpogJ8dLIO05jnmKojFYoX/sfbGL8Kf/DobZWuIM7gnKnp6oSQuDbKRg7sEJ8vhl8r0eyLzJ
LajUNdYrHzZKxzRrveGVm3hqYhFiaV5wtWPUX3UJk5NpSIoZp/4A9CzagDHuqJV9G0/dz8FpNIbp
x+4lwmbFMkjJAulv1EugYQ3eR3YZHMgxKiAuOqBiWB1NJRrGsOnk+nr53tAdUfb+x8s1b6diL4LK
McCT4bjC7Ra62j0kjPrLN0+0PA0RKR78w+CK/Sl7989h8NVTWuvhr+x/elAaJsrK31VYvTub/2nn
NelDvNIxNT2GeJYlVZZHXqPqnxY+TcAIQw7yHUCGAjHC1+3XOJ9o46c06SYeJBCbfo83qEMG0rkS
vKpjKzkqxOgXc+mSNBN/LBYfkZT8JOJ2X6TrhU8FJ2b/EHZEUzpb/f64wN2Ohuzpu3CFwHelbqmH
MSZFu9MZfPwoYMMwxLHNReYy1KHbjzg5APb7X6uXd2oii5yIgQgFy6o7xwCQJfxaCCfaxLq5hTFt
K5kHKsXEw08w5Y9r1Aqz6+Zum0eysPOFPvjqDAWuFNbP+6JD7A4DQzdjQvKSWJ51ZQs+cL+Z/bkS
oVrA6o92FhDXXjwQGluckSIVDv6JgWUDTb6uYqRq+jFwNRXmxj4iWMgDTmiPanxiS6nkf+xAk7l8
vYP5ar7KhIzzGWTB9H/YCxWQigFIf1FqDlb5n41LhyDCWOcW4YjJF8MzjmStF2WpFQl/HEVR/IA+
oE/tUrdVcW/9QKnNY4J1NPrD5Y5U3tqonaMuKeJ2FCtwRMmFMoY3HsMpOjj1xeQagXLaQMEIwTnP
KLsvXMX6JEStEYNnU0aBj5A0xKmY8519fCWI8VzDpy5VLZpOqfp7m5mLbqkqm8FYGDCS09CUf5Bw
avyAPbkCuVz1PQTUbBsnQmHtJO1k3N8V14R4XRqV/ruOWeEgYpUqo2+3IQkDj1TtPzQZJv0ggAE4
upb7PzOeYAdmAl+gGJAn4CNtUsImiIHXzNXax04NHnwQAtEhehRkRIpLoijdx+l+5SMC1ZHr0Vmc
O9XTlbViA52VF+K0jWAwL4ExDFWh+qRQeZL7oFc41nfZLDrLCTNqngAODWqwhNs/2JQL5KdZ2iBi
ZD+TcEel5Jkj0qJ5sb2saB/ZGpV6x71w9zPUY2bkq5uLslvJhfNWJfnDf5Y+2JfId0iPamzzd27Y
e42Ekeq4m1GOfbk4sy1Etwqnahq6HU1W8RxYGOrZLXDm9rq8Gcby+0MLxgpJetogDuiRMLw1xLvw
pZqj+L10TDpKxgUrwBqAz6+s1uiQTZahT6MKF4Nbo5PI/1+n2BI6xyww3jbu6CuZsYCuv9eUOvG5
PCSXAMmtkap+zza5Tg0SUfADChedARAefPCMvpU/UGB694a/xsLlXINMXP/ihSBpCBWHlp4Prbwh
Pr638g4Ay+kFsRpGBE5unnM3wLyTy8NLlPBkMZCTCrAbQ4AXcOr+8hdeRnceGfhM3hPo5XYdzvuZ
PzimRnDT/T/ESWwp1JSinWRzc643fF83LilwTJdbgXBb1R1GpA7i99uPhbZdWN2esQMlSGs/9Nud
5PSLLXEgDsZGGq4Nf6hRNBewJNaQqAS3vOa/FW5qULgnLANQRYIqI+w1J7of5Irw/q+Kxlq6jSj7
gQ6SJxUB2C5UgNWBcg9fsgQZZYdQwDMKA1IPRd0joHWbXUXUaxTYf+yibuJECnEC8VqV/YP2xzTG
51X2YtudM4bBZtw/db1cMqhlQd3P49gwY+8f6/Cv8vU7S9wUVm9I7YAwl5soK9USDTsw1EQVlcPu
k3BksxXvXMhNG1kLbVf8HVmoJAhCdwhI4xvAEe4tzigXezSpxf1UDjzm09mRdlrb6A1lU+9D7jfg
nYQ+gaNeQSBEdj61obl0wl5mB8+0AEfpzfaZAWrBiP41F6qp8bT6Mmj5z08lEwb1NZpzmHvb+U5M
OUwgKDaeVEnpyyM4KhZs2sUJjrL3eoThFirtZfNjOQ/UnEt8RiXKD1BeqfTLMqvUUmxVs8e+f8wG
D0gHFaQDsdoixSk6ESMh7/eP3OAF8DEINiQQ2q3DOCgphtrUEXiJMYJfukqqOe50ki1G8ogIN3hB
qer1ZCKbbuLzYdQ8yaIjLAy/NQphYN4tSvgnp9ut6A6xJdhTEPp6tqWs1TENjU+weN2/mCAvkjb4
Rc6SXvxKBibhd1mgbWC1ojJsvdtHhquLx9k/quRmH+UNNFJ4Azmc0QdAiU8irFisPfh9Xn2hcMZG
TTqWO+Awa0zM06juFqvM/zh6kt4+x0bP+fMfkCKrnQKeJLYKhKokzzzR16s7RNKs7CvbBAvUSSao
gI9PGbxW7MgwuP79Ub/RUEQg/+miarCb2pkc3JCObIMutmvnTyi2YbjCKW2QUTeV3xSLysANLulF
lvfmh0+ojGqNiuzc3znYmhnU7Dt6mDoYJhRVwl+oylOYDgMcqTqMEjHCAKwD4fK1TugiFfj0CaMd
lk47CbavDvu+JGAesFUzJZygzWO7x2FOypxBzTnakOpKlbucgg5sdaVPRRN1H6qzSsccQtOpLixy
bRpnZwwyBWqFfN4OikrnFgAK1R66qeMFA3/i0NoiekTsPHsPJ9/3ENlHz0I24DWTAjFPan9LzbJO
Sir3qW/+0bmjukatl5KU4AkbxR9QixYw65NvYTh4iuc6s9P4ve0HoXY0dJqm8ZBRuvN/ngGiYcjE
gdKCvXlyQ1BXwSQgm2uM/zFJOOxs06/isIExyftxL2mMp8E9O4EuF0/s9KZQCN1sqftv4RCkcg6O
NeAurwGZbhha8R7WURp+xQ+bc+j4pvHfAcdaFe2BPpeooo1TPvC1vAVvyKdUsv5ambnt3Bvk0Q3F
9V7C8eZHItB7Rz0L33ad/HdVgWVMjnTR5Y/G5eeTJW9gDKx1JNF3Fsm9J4nKc4kPrdX/jUJ7KI6T
6hd8xU+AzsDd2cKmXaF4UB+ngR1/DycN8o0a6/tHGYJc/+Kafm448iCn+1iRliaP/08IvZybH/U/
kS3gdW4TCNnrKF6U0/0u7RM7/7/erylFWWw8W4WzNUDD+z4z+sZU6KuU6fpxeyPWCwIUgGXtkYOk
m/+nZhRP3ZqLOjoDjZBUcJJ8/MLoqipIWL6PZe7c5jMEo5CxPP+8poRZPmsqZX5SrTw4cre3Gbeh
f/4uM1RuMjtjcaQ51afJfslRSD4GwwlQkhBS9atM9gse5pdsxCVe2tcUdWp/GA6yMEzDin++xzbO
ojgjlDC6sjpEAv5dpBUZ8x79r+b6PplY2Axd+8ji+JF7qTqhNAzX/ON9IJ0e7ZP9vxBiFh/QHsf4
aWPs0+mk3CwBCafIrfyaFQR+PMuyXitpNvEXHCs2+ywOc1ZD24KyAF5rsndokg9WWJLS1egE06EB
bxkyH2ADcU9RwP8qbX3Up1cD1O445Y0cxSXa4qaStIhOrFFdoAQT+4gNIkWF9t8T2DwLqG9+ebDp
clMy8vRD3hdvr+aJln3/DBOdnjooSfVG3rpIQtlzKwVbvEuwN713qv0Cdw9qMQTQQpOqVVrYb9WR
bVQNY0OW+bWp+SlNkUAncUcQ4GcpQ5NlWIrdaJ/J1IItvH3JNCTfx8JGHBDCIPCX5yT2jyP6J4zW
OXTadChg70gcoaWdoZ5psPvamx313oCMounuG4pKb9sTmyqxQp8nwZxt6auMb35p8PwXsTTnGj9G
2yqw1h6/9TEKfsIrSWgrE/TXrYjMrnsuRUDiqRW/jyresTmmaImGlfuCG39UVP9JFwA8c49LjL2+
pXB9vOVQ5S0vBrcrtVf23zpTuirdmGbP6CL1wwS/qqg25ofuDOuJwlZEKCLL/HSksMYJvSDWZrhx
4KQ/9hSzSALw1gm2RLvov2b9wBlz6Bjw0QWnYBrqmgUu8vSb0qoMcxQFLLesjw1vxhxzuYmU8QE9
1h4VU1lB39D7wUz2KPqDmnvRwFstNfswov1LlZfAxGn0PpMawW5774WODuXu9Svh/BVv0AvRllHZ
OMgOFwAg1qoO7R86Qy1Zq6zwH10l2q9aNo32MSgljL3nIBYO3LWC8YrEglDW12ntVDRdbBNNTojh
SiIN/6ifrc44X3LVP5q8s8aMA+MKgCXKcwYPo47ToFWr/rvUNIv/nPon/3L4GgdeQYvSMazO0XjI
u8Jn1TIxH9IeThFjP3WMxkhs5d2ztsOD/gQ0GXHZHuFSR7vkmCfd9eAeyHsyLP/iyZ0XeeWZfBjZ
GI8iPmdaxP35TXGht0gAHudFopKcIbQ4cazi6qauxN0GBD7OThy7HhYUMMuk4vYLw5taCnC8VwSZ
knSpPMrDHXYrvI33tlCvynUAqNSik2j52HQ3Oh5nfBpNz4q6zl0rvzfjZpj6t//O9xRYJ3cQNibC
y5Um2DROy4zlIgIzORrZ9yMRXHYr/99G8sbqz6QRH8gVzvJoAPXCjjC9ugoUkeDFlhbmnnyP5F9y
91hYC3aWr94WU6sUyc+YRrnGPjna6iH0TsUwz/DapxG3qywY2NcsVotrl86G0SGp7eHIg79YtAfP
l/3i0zuzsF3ntRL60I4hMQioxY+5RVI85D+OpkH5ijF3M885PiwTu93X7jH6/CeOEnzD1dVXZQoP
ZTR5Kwz1Pd1wEqwWoTbGEPnlRkwdVZ2JkxvaBpFRuMVlSbiFtH+ErlX+ZzIvWpcQLud2F96qndnE
3hCXkqIcOzv66kvgdLMfCq7SzciPN3KzkREXt69bJiQzN60n7E5WqjFsvVTNXOWFyD9BZy+fBt2q
liJM3QZ3qSGZVOsq8OwcL098o8bdFRmTrG1UdN/dlwaIxYmwuh+lY0zzzgngXVThhJWAh0zD8Xid
gtCb1Np/nI6YqkqJjMoMfAdG5oUWR9kHEy8UxtlSY7qf+H1HcrR9GluPzI+SjEiKSHidiaVz2DIM
Ja/wYqNXzr8JyjOuNLLeomqvHgpoedCuvuUMiRAoGn+YeJOk95He52DZ3fX82jEVyL48R16YFTp7
bdtOgU4J8BsR92KOfkQSdk5Hbp4RYA9uBHd3Lr9YYc/WEosJYVU6ItESmUIQDatRjCt5foMyACar
RQBAm3gZGef9Y1/uAch5Tiq+VeordzRLlfyUnYZWK7s+Zmy0gJgXnQhb/S6fEY2o+nY3RyvPeHg7
5NDiwurznMGgq8j+z2recoRY1Puy/9NFnDmoBEo/zBZ5UONT0+DkjIi45DiIb5lNT1yr46sBJ9/r
uVjWOPDbGLpUuZHMbipV8MPZZ++aj1jhpSJC13ssjiE78PXar12iAiHpKaUyXg5Kl1buLB9akoiT
ZkBfwq9emtTgsYiJJ9OrasgV30dxDWuFlrSCmk0+O6CN/0ScgcfsQw2Zoo0yRsycZBma9t1mD3RC
ShCDnu76E76m4YDxseh6VYpjEfudEx+RsgqcvNe+6KIKuBboWAhbHLcuS7UWIFa3sW89RfgNd8Fa
QFFCwjypFrev1dBTWmbqNpDVFFsJik6OG/XkY9OWF2XIAYDQ6GsbdEBUo8m4yW0KhxuGpcjj9IAv
wTtambLHmWKl+t+pV70vdmFbbX8uUqf8BLovKev55VQxXyKv1QQzjvhhkb/ORpgek7u97TTKF/lr
9sYyFxiySqQ0fuSOclrgcP3dRkSvt3yfAlMoc+SChZbV48MFzVWwBpp5W7GLH0Y/noR0tSquMTyo
aIH7KfZgo26lm6DyZEdshKnbgvGEChQ+xxjSeaTqI5gBGONbSsVGK6V9APofK2G8cM0MgGCWoZeF
rai8qtFqsMOHb6DomoxHWQNt2Ajl23AXxY7x9zH01GjE7uyJeitRDBSu7uhyLFwPfoiEgPjgl6cL
eQpx1a0e8t/8CoQB9d0kYL1JhJmzUkJpNPsoNTDAGr6EvTYTVSt8Djmc4NbssMtuMwaNsSkxpOEP
UYn2iHfEYBo4EXYtZ9MofzOH/NZNtQTV/Vr0lARZHDA0CpuUMLSjv3+kdxVPtsPYMByzYhxVWPSM
ZP0mMtpMnl+DzdIgo9V6rn7dqNkDy1/QjpSXSVD8m2/simCOfagIvCuWXfkw+SRU0oSd2rymnfk0
bAR0Z4/WqplU5gOkkf/F8Zb2tSCxCYqtkPgziZEysfaaLf6iHKav1FtfNgB5Ztroyf1NhpxOlgoG
ZVZbWHllZbK2rBNhSYxU3DG/t8FBDpp4pUdmnsde1o5V7KSmc7agrBW6vk1FzxULQVXGr0DBN/Gm
dfEWjlH/RmkAvLobkrL2MuDEfVfQUTuhcdIVV1v2+llZMBPDt5/af96oIujoflF+LCk445CWlxSq
ODy9JleL8VXnR/1FChQjME365EWfH887v4z2HuNbGmMvUU/M3EKWE2N/fQAjUkb+fKAAIH8IZcAI
2fyIloPAAtsmaBj0iT0wGJa/iePdhzwgRWMLLrP9gzeg9mIZ2ryIoLu8WL6hlG7oHWHUiDTgVsAA
E813nQJ9uDwZYqPBRbBhzMGk4SYrVeyo6hB8Egnnr1iS2FAgZ4JW8Ixj+BlQry39SpBO65GXSvNM
tX7tL5ZvQqoI4lknbwM5tVQ932Ze1aPcQxRwC3SU25R0OW5cv65YQCjGLBJkgdiVbm6+bRB9/pj6
NvhpuTqS0iwq19Okv4qO8/zXThO4ukBEw/CYcmu/EHPqjpZhUDRbWF6YCHQ8oHLvtpMvtQLr9KgM
/sPHChIFP6PF7BZSSyIXCqI8kTaenPnOKnYXOnRieNfN65QxS4uGWVwQ8gt4L+/4BEoX2AhKHS88
a0K2GDDZYy2GLWypSXGBhH29Qwrr1Qu1gT3mCJQ/pPtfRHcOjMA5yQ3CCHHdqu10n9TctK2gIvE2
2+dq61MlbRQdZf8c/e4znjElkp5i0AO0jeRuDkcQFN/zQEZKYnm+XbU2FEjjkSy+DXUBr1lN8Agy
re24/+etWakhLjQWB4AjrmBE5hWHV+lhuYzLs8old9l4RaI0XNs8kjU9EGISHqCLDeEKuCWchp+l
3RjmUpnnTrJpxwiAQ/hCwBPkZLIuQ99Ym1U6+PXNw6JOjq1PIS8X9xe0o79Nn0CixSAhyYSPHa28
/VwJ873u2WPEBMwD3/iqhG3EUO22lXxBT8vq0dtxjq+6XcvnQ4SZ95Jnb1WKDSPbLLVW24DAoYPc
GSknfaJmynC/rUX1ZdCo9MDVCzW+YUTRIxM27WmQgteeOvCHAvdjW2PjHpX8B6j5VZBEKq2VJSO9
Qoac7z2g1eQ0LZJD+nUH+OM04kDI4k9nnkeF7usvtrge6vzL1GfB5sQbnRC/ZYY9e1k9JR60ItLb
b/enrS6o6TbICoqRJerRd6YGHwOmRHLkuJO++6IPSFWdQrqut2BQq+cyFGyiI6w3LDmNFwYKQ/+Q
2mwilPIyx7kJ9dLdxI8SgJFqCWCYqMErzGS/WIImgDpwndSTP1ifWsrQAS/E2NNBVhJfJGLuq4nZ
K0bW98LZxJwyJ15/wGtNbm6VQQ9il4zfrrbnCkvIOlQeMnwd1M2j9xeqbuCojcM9j1MlTEA1XFXw
3T5b8KscFAC+G1ILa8e6OFXsfEAwiGLMqQsGlanvo13WJaYxgkNxn8E6KlsoV69ZN+y7rjLq3swd
N6NqH8x246PdopOCeEneJrW6YeTfXAcbeTqo0PjV/7kkgLcdBC+eE9DphRe7+NHGrZofL1ieefWm
Yt7GzIdRAhkT2Et0PQEIVgsJC4zMuDHkwKnzmmYT7/hPLccWbU7Cv3b36sBFawoFs39593D1dLkU
dKiA3m7o/apnAOjW/j7kXKP7fdMhJxEtVP4Y6LCVrwsAWPyHgLe5H0l5Hwuyd6W+lBW+zG+a1xeY
TY5PC3i5ykvRal5SsVawi7RwmgIE/IiUwIYkHi+D/0JY6xmlWXtZweBbZapZDzxnRk8cuyGw2iqF
RZc84nZWaYMJ/3SBoM+VQ6uDcfMGZ9MmWAaJhxJ6VgcSzWf7mFLXM4gCOeFy+B7GWlMt1riVC+vw
eNeaPr1TnJIyiTLat2mIDlT9HpfFURp/30rPuB+UzsqDXLyeh1fo+wRGcicchiTU5/ZBw7asyT4V
wym5tyipVTSfV+PeKUqqf5/41Igq2rLOtvrxRG37AYBqdoos8y7A7vA1u8Wexk7lHBuK0X9LTlNm
aenL2rtEHP+7P5sWdaUhmDe5bp55oRMgB+m6amEeY9tsEUdXG5h2zbinjgAtkjHHupjPuXjf/DUe
3jMAnFHfI/rrDq+3ynKsVUSfEdRsPgxbR/XYIjBS47QmXN4cDu5KZ1LNTG+l20WixeeMFWfoDhkI
EMZMY1zL7ROhTSKrCRraUyGGhtqdM7jXo73EYzqX29F4f2O45T07PssSSgzbVx8wV9fS+C7u5q0S
GMfjEleeke18LaLPuJmr8zh1pmYUzDO2u8dzZk0JgGccx4Thd7iMxDFwE9WkAEyjKT47Lu4pjKWe
Y0sJD/S12MDLTx3Lm7cXA43uy1JIkYMPnLH/6CNtgkSDXmbkxRtrs9ndDUOld/wEoh4JUNQe8G7Q
ngUGJOzidDlM+cUcw5icA1R0hEDGboJ/hBjFed66NXQcDR8nBFWbwU92VqoRKDLWwH2hBoGADFUL
GbfkjlegnV7ehmaWAwhNK0DZ7i2aVjNUEBO0inw7/saASS9xKvuHl0laPF03wNcx1BeTZlYW32FJ
v62Nex+nmf5ZMSwlnX7lf74VJtH5OmNt/GoM9lbPAyiamqhei9vpMAAK1EqmLiInvDfNvkCEt10N
osFrRIKiMFaGAW4mVKGOThin4AotNwpSHftt8OZzU7VLW6FKwhr8lFqdM3d/fRVswMdOD5LoA0jU
WgRoh9SqoN1AQu1AJTdiGlHh+ntsWU/4josly/RE9/av9NCBCYTpKI/y4/ldO4URuvb/PnoRNoNA
LAtyj/EQyprug3jCGbhqxtwfg3qQ1Y1aIYO1H/dhu5NyeN8Juxx5ZlNEFsh0jGRmHlfC1kFQT03z
35gdA3mz+K4DLCIQd2LMcidb12IkeTA9r+j6bo9lzS5fl7JqsVDdyupdLEojrlSAClEwakvuVY8H
/7PLBFWXeTDAuFGBpYUF7LDhnatR4F6i/fZMPZzhn6BDfQYGwsem4E3VBlq7VLuv6q2w47QyTzk0
ZApxsDwfGBeRUCNu/g/JKkCbea1OXmsMJgOcQjuxb7RLGfALLUqkBWe4qGeLO6A6o5MWJ4Icbl3d
cExQno6pB5gzNMPdND3io/zsxTeV8i6yKexpt1LyjLOgdnDW1GhwERnKA8R2w756OayJU/BMabsr
xCHuuuH105pqpsAOMijkxFueFrB8B2pFlu9klRP6++9SOug1+Ntgd1GNrlx57UaD989wiJX1/AMN
iK6HdmhL/p1BUWqvhKXd0ZQr8WATgnrCcvfCAjkCDbJNCcPc2wc7RqGIKdvMNaT2mpgWZC9+1JOJ
fFIr3V0KEr+USNt9PNLhiTXUzjY4gK4wOmiR1ldgTFQQtWvmZG3CA2tj6dmgoqqfkit9fozZmLH7
d87ockK6vlDb4GdfeAfFokOgXriwxnzlmNmFlKhROMAG8VToD485Bnap5oGeBwNHryMpKR2e26Ey
2AR//iGMf0vLNg4nbdYwwoO7VBUNAeBwk/NSKMurgHpaj3JatN66ziGuzMl5gvf7XYQAy1L4xP9r
qqOxCAQBi0F5dHCWJbvcU4BsxnoEqv+pfbvBOme8wBYoQQ7toi/q1I+yf+qCFuG1OZwWmZjp6zJb
7Sdn3U4cUBvbQXVda3pjkE73y2elS/EyIW9mgymXpG6goo/Kp2Kk183PQqRE0N5JTpY6DxWm8C6T
OJbcIyTtXNrCKpUbbREoxDQDl2/wowT4PiOVcUcfeILMzA+TJP/p24Iv7bkT3YS5uh8jx6ZdGdM2
iip4gFBErJAKzL0lW6xp1zWnRBIWSlcOJpoepK297Wpx35TrDClZf+Sl9opJcbGtDdOMHY8pHsXM
Ll0YQwwllD4NzMPAzTAtTvc4g7lVv51cT0uYTypG9TSXAfADgRd7KiUOWSaqG9+MR9KAMzK+zY9b
Us0DFdfDYchz4YKcRBLRDW0CgIBWoj4IL2QzRfOZodVbpFKaIv2nuBV2TBnGWf9SIHi4NLlnBhBs
L2BsHs9XTyJTF2MsDlizl9i28iD1ZK2ff+5uSXyAwKb7EDEvbN7nHuiP3xAISljeQp0sKFGqek/i
q2Cv4dgQ/dGsTHe1JLnda4zQKeCfWCSGSOyrTEOGl497ovmrNr1jOtFwWd6pLDFkhU5GONkPC98h
NA3v+BmB8l52nolJ303lOvct25z5ND68eIZ7u1bxlY5win8l31Cs01Hc3ozBvMqv+SZmMZZ4W+NO
ITSgK86VsRVwDnvERe+8wNH1zQeFZtAp/J4pxYq3Apumty6TXOtw47/trnisb0+DpsWJ1L4RZTZ1
JTzGzshkWp4WMKfL2I1TWQB7YWMfRY26q4vMIxf5gDJRBv2f/P/2Z/ILg0ZeGWk0dOguLScNb1ID
u6Z2fa4oFAeJexsU5DAJ1u63KMa4VbyetuD5KGjd4IkLdRvMftW8bwzMsXUn7cObd0OzwvcHfydi
+p/IkNMW78vOAkirAWkcFXrojBiU88djPUPSJlfSxbzA0xbhMGJqT556SKR0FShM1Rx+kcIRpneh
2neK45XBmNd4m/wusavsbeCwwv3bZHZct1MdRH77EPNHpxHV+NSRt77TOvoTIec6CRyGj0I42x+d
Z2a5IEPMJdsdlNpQsBoPKCW65RI+TXAi9xV1JWy/7q0vwVwFgMimzzzGLATHYiOCmNK64/ur+Hqx
tcbVKMIlPjCDsoWu6SlRaxkQ3XKtOT75v0TOu/oputC+Y3CI0eg3o5vWfuq71NyTwT3iNmeWLxFR
5LOPri4blFtJCwWGQNgCLtPUBceLOrvQ/t4b//KrJf7esSzXHMUNw9Gu6P0SypNqlAUZCXTwq4eA
9ilMHqaHy7RAlAkwwl7ivVdT+q9+uFiWBn56/N0W3DZhgMxRJuPzF2VhT8FuorwUzK4pmVn5DLJs
ya7XmyjXoVgbzEUnX7GprCyKAZdbyOFuruNgfJwawnzWZgEveipNE6SIPFouO7SC1SJQy2u//WB9
b7QqesTvJeCTvP2esERVv7Ow43h4xl17VT0Wu5cHixWA6MNKR2vXsus5ZrlyEjDPusojtZB4CWal
K6K5vQfOFLQQ5ANPczPywo5CL3AboT9P96HVreu5BE8dLzyEauTQLOv2aX0LqBJ98zRChVB1dzU2
CikZU7+XmSXoZZyJTJnfWpsrjX4/wmBikfTJQEzqAhmmqe6GQhgzLMvPLjdAXsf8Z7o1XM4A1GpQ
xhwN7CmWOFN7E5NGFVEggSqNkCyZ5+Nzd2nyaUNO9f0gykRFbdXGrk3jRJ0VSUqcejzB2PUUD6qS
k17f7jYwECnDVpCMMmXWEmzByZtK1X+u46D0C3VNl8cE1NgP1Jr6Iw1a6qVKOpN2733hH2fNQVCl
bMnjCDDx2O347wOE0wpSubjcgfb58VExBAsazxASV0ZGaRTgGpCEW3u/vSr0doAteLurw2jCIkC4
Tiucgs3AKa+RXcKl49GtMoEY7ZrOi8a4a0dBOroG2zzrhFxwQm84hp+7NpwhB26aJKgfvoV/Wj6H
eaPADEdfs6EyVs2T8ivSqKA6/juzB49KBV8ZNgT1Ny2olU6Xugxgdm5jVdik886A7T++8KDNKzGp
l25P7CtZz8oZO1nChZamrYjqTfRO9uauY0kbj4n3lIj9GD2zonKD+v+FdJro7j2n1FqxMGExzZRV
Nu7i5/TVrKDrsJf14zueXFoIGNTTUHsV0YY/m1nzlIs+LBZCkRAAM2x/5BG2L8Gt9Ug0GsWNG7+Q
dEFE7XupviiAPsX7ZDGeF+UgwJktWTc0WYAWX7NIM+T7mXwXVrlvhhI4rnOgV8cREze/bhlwc+he
CboT97+LdREsrZMQMaXOoYiotDHeARmsDUVHSaploB2zQxWTeyyyu/PtyRUKpoKb2TMVubL7MfqJ
r5Mb0BUUn97iDMTt05IAljMQyKKnxcBIPxMWJARu96qg/WlcQMirGJEfVRkAVFjFhzTPLtzS4VQH
qgaWuC3px+ZGKcyG0cMQ9rqfGO+94Vq3c9Cr4dUQTv6zfCxWUGccHrCGb1jsiYzONY6fUjSpNmJH
SBaAJFs5hKS21roNKY9ivVwWUx40wXk7Xh50C6oJdfLH8oGoeLuoJXbQxfXcQB4uFBjeMbGKEGEE
qjgTeEGwWqqVTHBVPUF0WjjhKHqZGYI9HQxSJn5HKhnhemVpoO5UB7Ld2MexxgBSZwmIQ7v6m+BD
jEF2x67QTcYKV70Nx1b+tXFsjmqKYlNduggz2Pm+9lXvzu0DjrAze6hJ1DDX40qu+Ps5+C1o22ye
yj7AdeltzKYcW+jUEtmVNyIlepjVhFYntPdJa3tsvXlFUmR9wYYtMp/eYAJhCYmQbBfVMkdXE2Ls
OwKJgP5xVsHrAD9nUBExDAZJL+ONuy/irEyTN//HGVVXYrcPufXvc2tH4lDOM+Wjt8OprrQYalO1
nDr7lSqKfBTW9XelelMYf+DDJCOtrZ0o1fyyT2MwwxQLfwF+8AEGp6LXZJbp3i4SDRu5IB2qs0qj
+/HFn8EmZCnG1nmEuU6SLSA8nb5/gj/YYmbHRkqsVmDkXFb6/m5opyTXXKtEY/BKYhecxjrL2B2r
X5hemaJEyE5afjdvlJaykpPbHKJmAdT7B6AbNJyjgwJjRy4Uc7hH8N9ZzXmLEkvim1TZvmbTdaoD
4s/l9uyA4zS36NraiUCMYoXD1RMnSx6eadsiBPv2AR8vHPkkWoPMIY3jiNAW+kEjJGb8Il5/r7pS
3r57Q70Xw/06+z04bfI5zIx6P6iwUKqCouBQy6fxej5+5hJrm9++IRHBm9qrRHAHlZ2C4TeO5xj+
avxVF3l6nlGdSpeADbXlPDgmCZwfsPoMJBhADyLe7AKeAWg3x9dLyp+y9o4gjV4dqW3lJFhYspbj
SR2c8QbdZ4sf4jyz6jglfF5pkHmel7RJJB3BQAHxmNekb3Pdh77kx/tjNJBVu6YSUjCcuBp7FzNH
jdooa3rBKD8npbBDHo5ujRfznfw3QzxTamUbjpdT+eZ5rxDlUlrQmVeMz0MbAJfrQ6Tq4e70xH6h
VRVIZOhNPgytHpqS3NoLz0CrensvWM4X+LS/K2JJZ9NPEcUUQm8tsxFk4WptFnBvmqh1q3oOZmqD
nnscWAVHkDRIxQ2rbwh4HkhdrEX18MIfBDk0dctDIt2B3Stk6Az8k+LID+5R8HU2P3e8mbXBheZR
9/3gClU3320IUuBQBgmqMfh5ij7OQmH5c0WRmuMUh1osonGSDKfR+U/+R+L6PbZqgNVyYL46JT8m
E6SpHY3j4fe27LSjS/EGTtSLVhso2JN0EVg1/EvyDjNTSg5SLUS2snp39pboboznjl9F+g8BAuHs
BwKHt9pT/22yBuS+qCKbpGeC/1Fu3NWI92oaSHmfWBBOuf2RnqfkNMp+KXbTUrmusWJyvXqaKhb8
LSqF7JZfKCWxAHj5/e0pelegDHsZ/yrdVbZrZISYo0fLZLedFqQwaTSLIq/rTk4n45u5UJBR+4xy
TUb9BF8EQge60XYowqGOqoUf68fS+/5BqRzE5eESlIz5aWPyChM1TIf64Hr+9mW3MdwCq79qFAfk
LTnMpg+tHNOsTkskbqbDSsxZKxpJJQrwpL3oXv1uYFY+eBc3PdjUIN5gMoW+yPeAvHls0DkNTFLq
W1/MYCjYd/6jZce8MCWM06r0TqtRlv3pr4NjgIMIA2sBMxrRRcjh0BpiCfGRIxgffHm0LBPvkOhE
BEv7ef4bvu8Aw1lo52VWvs6nMjoKEjbKYjafuxYXKr9trvUtQ2zFWumBICiz8sNUTfLDeNAT8IZT
hk4vYynOWd8szHH7Kh0ayBx1RlG3+78PYICIQ0G4u37Ldpx+5nuoeViXW/s31QPWDdL9bIdMPEhW
6x7YsltTAsD8h6POZOgoJ6VHuERDp7x4ol8SZ2iqznPdiS1Og7TsUCY89k2SKqqB0GwPYW4Yj3ak
yqObYCysmwU9FZi6qJppZfGJQrAQouidFFhsMMgJiOjBvjolY5Nfzcu63fSAWJqhLCYhpZXA3Hv9
HkU1ZAB3xRcXtl2uNq42cawBvtsnQ6x19PZ4dUnETSu338kfAllr2z+/F408UhFAHnspS+KLe9u/
HtE5o5Noes8whGJFRZUoJZ8bTy8PKRNb9KFWdsmN+Sk1Q/COZjUCcsPdxKQiteESgE13uZlcZ7lb
IzNOtVUu3QT5rCdvwnCaWoHwn/4KWgNB6cstoG92x9oZ2nE9N6wxuTY3M/RSykKhnFldaBysyDIh
jX5/Sgltm252RrmNn7Q0TsLbUNFXpa3DgcPkRDGEim745fLqXg99WMI790+jTO5QZJY1QERZeA19
wsOCDa7a9jPfoDmXQxDoy04m8SWLx1DmeijM5mz2I6FyrBT7s1TOlPV7wgLHIO/v4F6sqgz6ddpB
2FcgZthJmOblA+vyw9kmsrRdQT5qSBcNKCWkrwPdHQFoiRbiIxjJtu2FXc8P2fsNPsEsPf3Eiwhx
frh0Odc8UnS1eXWWooxhV/8s6aWYOpDModfVvcKGw84WS3I9X7+cUW4SZwe0TDPnX34AVCF+ax8r
qe4JF2HqR4PZlpwzy8TZb4+/04MeYJGqpyBL/de8/NIC9ogP6gZFmnfSBxRF25DY3Ptiw0gW8QAg
pdGkMfjIjffxGkD6iGexlNUZbtjd33ayi5cphpsytb+HvoNl1jj3s9JCrR0CANJU6gu/kyjZxr4m
6YtSWxNyFaYeVTCE337gkjxYuOXJiQ7iiFNOw3825JIpHWHXvx6oQJYZn1ef+hIuB4JFY7A7Fsoq
MMzOhvB/IBZ9SxeFOzpBH3+HntBXDJkfnftx95MvOCmKVKufYJnAazWRsHZmuU+ZHrxSUZyAMwSD
Ll0MA3DtXL6KfuiFflAZAs/djR3OxDk1W5u9Tonkdu0LaY27et6NhFtW7TYWR9+kqB2AbSe8G168
MicA2cHkP3ars1u1wk6YHUJJDyL6XGZpYRDwwmv1OaPXm3wAfXvDut1k9RG3o2CQ6Nmer/rosSFg
gRqGsOcCQaLfCHIRn9uU6GwoZ+X58UlVebyjiQZr4qEoTLWov40naoRn6FjqXRHpVQBnqypbWbaM
bGGZGhZJ5LhXHB0hSLvKZLQhTGd9VcbWwVvzacagEJqTjwJAI/GFTZRK1LBoxhRozjSSY5vpojjc
2u+2VH3ETAA3J1QpOFsLn3iKmQX9U/YFTciihgphloSebsafnK3XDSImAczopEdFG7L+9GlQKo4j
o8BT+yX9Lb1A76wAfJHPhyWOGNNJUcK6ddmD+pBo2TqpZh4Yb+hJEdZ6eYjCJ4gDRjJeS+g32+lP
Rt7is4E1Nf2Y4i0hQrFJPlEwEAxWzJXh5zYggkNrU1s7XqrnWPWEBiYYIsSkqwVWXH6iKQ5NS2ER
zUZXawgquUJL9PNQi2ElW2QjvO6cdwDNzxK+luG3kBU2GPsyoM2p8H94uBM87xdYsfu4LvRrYwlT
1fB2B8bAXQCnyrks1HUMgIvBDhz4ehIUpliRlGEc+HuInlP/gxh12aIwE8huQ8onhSY5JxrHn4Qj
G4fLf6hn7h2WIng7c/2YEBigPUw5DRxhpxdmwF97NYN0T243cONq4zru/XNUJ4NmIr/xu9JTrvHF
7QRQYwF+c4PWrHUFP8QI3+sYdgAaCqRB1Py3s3uk5mEQXta5l1BDbixRNvhfep+Od2xabv+7GCI/
H+8SQ9oitvA25dFS85+di63g9CYNq3y/oYEq/P6TSrmUVQK9ITOFg96IR7utpzIY0XxgpTdqlQ0o
UWm1CKKTXtXHJlgQtP5LFk4dws1KppVQqXZbD7Nm0PSWRdA4sNZNbTMoE9uZe4BZjEggygyMpYH1
JW0pRnInXUlE7FQfo5hmcI60BDo8sPhDIELEa3DT7V7F5Jg0IBYGm7ZSHMxq5wI52d8MeBlXxW8D
+9xfQzUJsZBPlvtdi7MyU13Jt1Bf2LQKs8XiMhbMJZSgpl9BkCFRKKBhLdgNc7+9/DivJSkyfbCy
izS/wnSMD5BKk2k7Nt2f2M+RqMDF/Q+PA++JML3yqGG5oZys6W37u/FpcnvFbI0RtLr7y12WyIJ8
GX9J/kuJiy05pvXhbfM6EH/81tYzfYoTjCHdsh2wTI8eZMDz+DDhzH56SV88E92QK0rCABcBj7lo
Y1zD3DG4bFfLK6VqBmDQbg1cfz/eBHb4LETXvx5kPABcY7s78zYy7u9IzwVQp3sJ0IQLyCKlWdYq
PPSPyMOIrbOfx9fZxzCNk+uGTEwWhh7FHFJMfTTRqAULHuAtLh+genK5ubxRY4UnTlYxwub4cSu4
GU8L1dFRaV8f8zwyN/NYK+nXvDguQz8lIt6KLwUXSXZuROND3nWRBh1R2ruMOgk0NOQh2jR6y2o8
eTndC6b3f0JeFB+bsPLwZGDosPvPS/AyK0Py1GmRLp4IiX2+nEEpyM0MHIHUounLMQRF0YDbTPjb
/87xUsfaM3pGctDPCkFNEHUILnFWQ5M64oQ/Jf+BGDWsf+RFPFUZJVPJC5I5r7S5Nbx2k4Ojilwg
0iu5ZJvrJgd+IxNocIJxA+ZHzE42ui/phbfo5qJ5NYbRYC7ewX8iugcF6AJlvIjTfucPYtfU5G0s
exq9hP5bOexeuqqcU0qTLzIleDc07l1Cqjxu7H174auP53x8UDthxilvCzBKbNwdh/epAiwZlK4u
dcZlhKqDfzK0hUHXij8211whTYzzuJ+DgkntbvaeQZ3bs7BevOBTWFiT23Yj96yR3L49yrxgic0d
Cu5dkDfkttCRrGE9GBm2BFLIRrbnOFJYFtC3CwbdoW9IkIJmTMCLw6Yz2pKR+nIXW+LTMsH+JVc8
JQZaU6aIqGNqIhyLnxeunmtWFTMnPc8/J3VnzjfjcANFlh8nlQdUTqHugasIfs3yfPKgjD72SsIH
ih4M5TTWJvMELVXdAaDkl477JQPRz5S7uiQffRwCSHZi/vxmt69GggkxuSAAA0JNHh1uyaIhey14
K829mRO+d9eLhyHrKKWoyUUPT+cBL9Fn3qtn1A27k/oxcnYfO1Rzepsx/38sCHa8dekRbfMqNedR
NwDLKApTvc5LGiyUs0Mf+i9TzfWF54pmCvCKpZlSK2aVA9SBydK+FPjgcCZ6FwIPiQVXlZTiKAH1
P8Aesj9l1ncmJb8GIk3JzK0uoeI3uVkgd5aY0zZdJx9GK/U+ThUUnxvr5qt2F/jakS/RjiboySJt
B/vJdUdvEWhlv9yiK25ODhUP4CZGgM56n5gfeFwr0TxukpHivooZbkbPzwqoQEh02rzCHK+1euJ1
8c2pIml9hQLRkYohrtXbHUgZJzpXePlj2EWviS+WUWC58IEIoEeWsqIomPX/wH4bz41CAdKSpkOb
81jngYSxHDfKLqLkO54PkpRZ6bicSSgh05ygv7olyFbEp5zb84sdnqlsfOEq4kbzSdkg1OJEj1Fb
6G1xvgXCbslqW3Yor2JoYWtNgjHBm/B6dJSwZJOFUqNGOpApi7vaW7D+dYtJoEOcmYHVE469jFht
0vf5t4334vhBqhqo6q5d0KjpqaKKgS6gIqE4EtJeFmFb58Uk4YUPXCjOQbX9BEVjRzxHyN1LKaP1
WjiBnJyK+nHPb2o5vC6hNNeHDZ81UYQ9nb7axNPKzdo6JwuMHCVWTofrvkqJFbXjJdd5wlfOsxNY
3DDnPXmPyKqTKx+91AxAraATYGMVnjBhKGa3HJEw1PbqiVxnAYx9mgy9G0JEz4FNVpLL+5RDmS1O
DJksrC7GLKoTbxeMCOL+IsFZUUTp1sLmh3Iidf9xG+frFLJIlb3iBHcd06jvaspVdvqlL8E00UEp
vBYz62lqr3fbdF4wISwlu2dYinQ/N9mFuadcxrPeAeO1l2vpktQ7KjXYR/a1lBuEQUQ7DYoOS+iL
H5LQAYDXS6MoGTdKR/jhRYoGfLiGymB5qhKrgSGTrcolbM9bIBjUcVq81Hvl+pp8rTc/UGU+OSBL
D5ZZiZbe6iPmn2NVCfHOCciZuDG7zCWhE5aH8QaKks1eG/gwRUlHBpiRIBlhDvG1addoh4bhYNFt
Ar96azidNAogiHE3teA2bdlM0zuBys40hNW/EiXwcQTSAUJPAJmDifj+LtOn3tCLpLiTg3IJxJF2
eWRCVXTxZ6UbFfbAHE6u8luHZdDTe4wxZW1kfe1uCzUUhGum6yusjW2x/CqfdGeIRDAr3plYKnvx
kx8Cf6bul1zd13q3ykXghuAhPvSdAk72gU+0UC3RunJjNd5iwl56YVVsmlGa1i6A3C0JCTCDzqkC
GOZOIGUc5RIduRv7BoplJDbbDJZZ9NukgfD9xclIJSKFTcL5tg+tYEamzrNBwhvILQ3Ejzs5Khn7
jAOWNrcLNehxffArnea5rHwPbHikNxiR/uZwWoH9olEWufMdcWTTd6u8v2yX16/vihNpYaR5R1Ez
Mknvvi1IihqJ3RHo+2s2r9btjO+8VMo9RvifP/MVT9k+r39PRWZHyRlhArUre5a1YE0M3Z8ZfZru
7ZotKla3+KPsDTnF7qVr5VbMKgPOxfn7GUKqYM20fbKlhIRtI5OXMYqstbRTbtsX/asVwymYmuzW
KL91frZnInSSJW5GZm/LJ/fRbEBQUH8J9QpPMT+a5oqH9zcXvyM2Y2MKHwjS20df+4pHZ8GHlMBR
q0DA+cDWJLdskbcxow5Ya3vOJmBxOJSj4V8seEtIYjAzVsByCbyMccz+/A63PToqVwGxjsNhQCOt
GUwQB9ZAtCakFoRQW/z3m9vZbQrjLAb9+1Q1iK9q2JrWJhwVOqq/woZ9alm+kHZmCGD9TYIvP9og
oxWLlw22GL9HNP3QtRa0oVijuKFWW/T6KoK6Il6GlJr7v6fS+MiT3JIH+KZ6RMps0qrdDGe/EntC
nE9yymf+Tmr0cNvU5h+z0RwbykDYHSeaRHQ0F78T9jeFsAQSdZYxwYKou7t7GqZPVsfV+FIRGrrw
2cw8no1XLNzxgbjV63y+GBQeE6rcKVuyOE5wxYPohCl/erYO9+A5CPaplyKujxk/aBQHyRgEd4iG
HVZRw3/GN1qNXJ9XkyxLGbB323GsrZZz7290zFB0xTqWu0dRUT5gUKOEssF3CQFQx/lma1543n4N
oJIPVxrhLDIudTuMXJ9PoRGoZl+yZq8VAjatFYgV7fQPr/ohOBSHE4fZy50QTKVGl1nGvooHhJQ4
AZsEi0qJ0107tKSOoj3K/pQ/rSIQCNY+nmMbuV9VPrgfOyGp4Mp8tY/+dC6vc90OHQELzdnBssTe
M6mvtSdSLHYV346AbL7y3pvOfccHKRhlZENWHTRe27tGSow+0I+Kmc5HySgwDl8c3b15NiNk1K0Q
0OFCSQ0pmgy/d4RISSk5Q+aazdO1fsp1hIbEGvb03/p7m4nweeJCe9dK67BMJ4fYbElH2nN/rmJK
/Ejg5FvO040ygYp8fD/k9tvQ03EZOBO6oPfqtPI6LUN4YAkNLsuPpNJ5YZl1c+7RIy80s0Vu9vn2
0ylGWimuisfZZ7y7m6GzAxLGu3mWlydzhbuF0pmcAvfe/cNQw+f6uc2vq0SfWrmJLN4LZGsoeGm9
Mb4RYzTpuVDKuNSUsMCf3T3tXbTv+kMXCy/mvEYyPVcNVxhswZE4H300+oJ/PqfWODvJmO6u0IxR
8PO0u8V3sh3ECdeagIN7mOC8r3QJDpm21I7pX4tZWXbA2CRX87ZLMINa5ilP94Thha3ZVeanPxxF
FX/xVpcF33+wviaCTgGuShncvqjZqteXIFaN+uTrPK3KxBzbdBH1biK5SLXdobucCVWoHDFNIaiv
FhSxORGcOhFY1z56nuzIdl/3XGCR2CxbFiivK2eEtB3Ss1/xke1DvVciMzRu8PebXkHap2jDGANr
Jod3t6i/owW32nPp2CCoQGgBnW66m3pUz1uBYEnlTnBVCTwP0kwBmDVEMvSt+meRN6DLJ8vBdb2/
v82+yVeW6hsYEvDINF3RokcyqFK7HeiDx3TrTVwHAy6oc0R3UNlXCU6O5gKhQ/h4iPWc40D/LbTd
k3HOxUMe2RnzHr4lv3acJt6FFaVm2bLZdgP1dce/3755HCmmWLSFda0md2S1TZEl2L0XCEF+7zaN
kA7GHUr56wxm41IkCYQ25VKSfd3q4Mi3qaEZ9WWop+EWXvpgXVrN6DVw4SHg7hUYLx1ip6HkaOcu
Y/6V9qd8ZXYD/fgbbt+sWLfwHX2VsZF9qEmg8rhDZmnPFqLwzaPX0g/yqNzLgQR+wrlWu7u7c0pK
qfs1X1frguU8SS9cPKnaSinU4XsaY5d03LoSnVX1hUcYQLZFh6BoJKM75faYO9A0nCNV1zM5vDJK
i6svWxmyNC9gzC6lznE9Zz1CXIJSMhnYqPCnD+H7xHnZ/zPY8IWI/dCgqP6dkEsiiEfUTBaKDKpm
XySLVfkAmudoeRWEcqBshnKjrWdDlafaaoTRot7igh+j1sZ5VRAaA/RMC/Rv6V+zHeVdOcga4O36
mdbS9PCa9Ulk5I0aw/howUyfb0dRuwDM6/wpVhqIiHya2VuJYk/D3vd6FpW98rXzEtXC7Qg/ACU7
V8N/FGHyhyBN5xlmX3lYadj94V1AAa8K52KjFfooPD3bl5Ao1KS70bQSxmd7jNUp8vgRJuPeBS2J
citfSv70jXRJ8v1RWeALYyOsXr2ZzfAO0QmtzgI23oAZjrbtU4JnDgBpVVpgaE7kpL8rYkjMfuun
bUg0Wu/gefyjtQf1BWg4SBvqzS6nuruP3jzApuXroPe7wBSkJ/WTkLU67h2Z3jadWk89mn+gvzk+
BrpX7tIyiZvKyjT+ff+RYmAr1P9EZcADw24Pe904dBTcBqRFCCpr+XnkKYUOED0kPPDbN837o3Ba
ngwkqj7CTgRgF0mmY+A9CjC/3v9MUt00BT2Zrd0Dh9sU7yk/424Sa+hqG7vPxZT8Ro6nXAB+vG3S
V8JrSdMdt4nqQ83e1eAkdHhwhO+ZjlIhJGbVhi8sZdkWv5HPrOzFZmHEwtBNM/tTHVyJKuemlAle
+D7zcf8b9EaPVeyMd/0c6anqK7TX2yXMiPot5Q3f9Bxi2wAAZDBzXSSfKVPRs4SU8macC++DS3fK
jDv9pkYHm/oOXWOdXJg5GhgdfxOA/8TG3z8ztcnQvYpdmhxSSExQSSnKDgan/saGvq40mpuaRlUj
EbYrQgV7TY5uY80Lg08gSrtlqDUD6JHCHLufMt7ZfEPKlxup2cwrNqkYUxjvLlt1TaneVc1sXNRF
Js+C5lxXz5tEZGLJnAa8yblpqnNZeMI+o0b90gs80rL5AVj1w6DowtAoeXwK2kNZBYgn+BSgbIUz
dIelzXAesBti9yO5pI1FbxdoWnWkB9hCUIWOJ7b9EJ/rxKtK5sepY7EeYIE13JDYTcuvq3/d4vXn
6/Ro2ohaGF1WLBIqolIb7btewCJ+P4U4wG5EsvQwVhBrF1w67wH4il0eA8UCCEF4hAE9baxkK06l
a0uT7sQrlLj69WYDOxxciav5ybHpWHqxmCplGj1BrmfO75L+62Xt91ApHwmP4udeHHMmioCsJJPZ
dTzEglUC95AhnlBkPoDDcvmxR5Jw/2RsVY7FcP7uBJNW6tzZn45jB4ySkrImlShBLIFeZOH4HBbh
T46m0KVxlfr4MGyKJeP5uRRjbp5EzXK+0m7idGOevbMNWgNARsTc21oH1D8I0cXIRS3XgFqaCvvN
tsijkenc7EFhP1Xfrv23r2qdXZHARHMjZb+2XqJKE28ig+VXl6Lb1HCNmcj9nECVv3ao+ssVl+Np
4wT60nP9iLV2jsHCMLJIHUwU7XXorKS8eY3G0VxVmL9pIuNF7H/s2Hoa7/OchdP94Wf50A30QMgl
2ufox9YVmIP8ad/UOJ1tb5R7or8IM50lMmb2ls8d3SHXM0+fcFMBaCTPWQ3G4Jt/1ESTSYNwliOp
0cb+IWGANeo/oYQRdlQOTJ0B7/0CzU4kXRoHQeITw/+CfKKB6YTH57ZW8VIjvLGdHFZQAHfj3W9N
gRHpgDiAxij7jKC7tXxg8o4mIGKvM4IYjCKNf+YS1yAQpeKfSPQhR9gcC0hsOEdPf4M7++v5J1Xd
Tv0v4Omj7T3W+bgLbBoGUG+DlqBmibHXv7Dp+hJSKMYNq/Jn/FDgjio/ODC+JuVSWwjYzLXCwYsV
xSxtgeZOY91TklM2PhLPrJyqXjP3IBdp6Ma6p+3pSMNAUNFf/jcdRMKoHMTpUdqpvOdRDuIpE4GR
u5fTKMs5VdB8olUJVc/My1OFHWDTNnazrul5IqP9uVef6MPsapSa1Ntoms2ZuWcItY/A+ZYNa+jD
owRky0w4epAVTZLZD9pHTY00MBPVlzP1TEjsCLMSQvSgeXSW4VMTSoA3X2rULO7ZUm+l/twO0kBG
XdeuTsXIoE1KOJQhI2oB/BjiiOWWcHwQsF9UR9KIoN9eODBTO9HdoHbTBXBukDnZBmJIELfV8bgJ
zfVqODpuP2hayyJlXBqMaEOtSMrRy+Dup8QoZBT0ARBiLsmRs0GbhhoNIcLQ7LQeQ0MQezQKnLCZ
6i5MuDPL5umXgn0JuBj4x0Jglx9moWCSHmQ7xFJ5Dqqo02rD9dhuqmXgkx2m/nV0E6TjuszWC4Nf
ERMTJUNSqKRlt7IDuaiFSPApPfFfSxt5EAeaevP81V19o7TqCu9XxYKTKCyG0jC+ubbUmyJUqJLO
AbQXfOvg+tCUC7MGZy0puf9q9e1NjbFkVXkAIehID8o3yOErCZHpRUl3/M8tYdqCI137dIP/beSl
/PAqpAA6qr0Tm3mE3li1Pibnh3bvvi9v+hAmhnJcfNN9yeq1pWtkcWmBaQXstxs4QKRkMnI+0iBF
B/dFW2yu0Qc2vQcszCmJ3PgTYt04mdvB7MI1mn+p2bJeU5Kkily7jXa5ae3hjjfE1JULCpG3pVHZ
CEBGoVeFmizKWlYgcOVms/QvKcvh/q5hmVQ0843NgASr0LgiTNtP87qD7t91y66QMQ4tVyKiqM+5
0lv9JBy7oFJfDO1cGOoClmAC8EXFafS0sTYJ0tziU9tSiOL/SQ27rLAr091+UYN2W5+mjmIEMfdZ
iIQEvOavEwOAI5nEWcAhqxkYEgEwtmBvGxRNHB8NuxWeZR31Cby0DlhmMt+3b5/ZBSc2ovXzBhie
0Ov4+TjwW2Ani/rAZ1wfa4inr0AR8S85LitA0J3GCDcyNIEtQJDJGIDki8HiWy8n25AxrgfcTNCW
nJF1V57DYO+oBd2Qu4kSan2l4Av5g1q1AI8U0sWQG9YzNOLx5bPA3Go+44KPho678sKLAzX0YneW
dWYaMqj9Ao//WeuwCW2oNBlTy8eJxhnIOwNFaOh0R9YVWyiKz4vBj5/MowinOuU5rBXVobAbcpNT
K1vyM6e4jfdq01Kzlte+koptMM2pwsmu7JGMheWw2XF5fY4PSi6iFF5a+fiUuQqvsIw7NbIQpjDO
NZUjN+rAdR8p01drjsjC6vYYIIoE8kHuLq+EZoyUL2sPhdwDQ5PPv+K2acnIqHay6hEXIU/VNzjD
k1hq+sykzOgqn+hZ+CE+N76+rQ3RYe+/ZNEUVzwikL4gq96BqurjUlD5qOlQJspvGkjAz38ivFBq
fY8X731oJcjaoAc+Be5sZ6qZ8XBG1DZO6Ru22jT9oJ9GLpytswcjD+AQzm0uI7HAZVKPJnpxQswj
1zD8vKs2KmqQUxI2qELKC5YIFA34JdtDXHw63sbDqpwvjSfUGG4Ti429oKOhqIqzZLfxS+8EBuuE
xw/ENQ7aedExyKOvxs1DXJ3bgCzXhc3SVjGiF++6w3G614NjD2e3XNxBHJcDsmhZJ779rNLOIKIW
B/gGEIbuYgX1wdknugRaRYHfUwcny8RnhtBZSeIp5qrsgPRtub3voa+PSuykuXfV7vinA3ss9br2
S4zkTcHFg70bG/i0Y6Fg6bgtQE7gu5F6dusxLC6UBi1a3WIB5FZeLgp81hFHsk/EsMKwVUnB/lXx
8ex9o0vGbDrVTBPwgJFJAO8one0VxELWqS8HqPrEMjqyLHQkncOy2N3dvI3cJfJt1TowcIhXwm9J
KT8/mQfxq/l9EyctvjWEkGE0F1dXpKoCNIVlnO2RqDnFM3qCeq4VQ21ZlHmx7GPUYyTraX3ZZ/99
Ophy15poVC9ruyPEc40SI7THk1fE3YtBZt8sYfBFi93wwendqOtWWOVNT28HWo8r8hm90W6ddJNM
bhE2Fq5h/Y5LdYZqF1M0dwHxVmSVb+l0/xRIrlM2Wp97Xt2QEAIP/GMr780eowZFi5qnhL3HbHrU
MgALYB2LNzu3/SjVDPc9FM8vXDdY2Qvu0FPzRv+9nB8s5IEFCMC0vJn2AuGK+WfdpSHEo1CjF3Lm
rd7JVcQ9U8G/mlxDva3YSnGzBJhbAK+0+wE2gJouEwkX1TjDOzpDt8pa3LYk8uYZv18nwKf8fUu5
1xiLJuvUBQFqGaqrac5QIE1Ax7OBhWDTzgniBFPy2OXRCxQsGejpCHIHxfHW4RQyWEu40uwNmhtd
g6Ja63umZee2OROL0BF5UHuyXnaxUut7eJKfeBSd4o//CJS5ayMYU/dCOHw1ZUprg7oiwjjiVIn3
06zPAagel2xbDIjknHomMh5G5pFaOcWzXW9oPVqGBaIFDeL3J0qzrAeeuYLHWECcZKeiuvkfyL9f
oerpL+xtGcKDWuEruPeiO4f38wqfcYMskAKUx/vOaIzJhDlgAQfryPqA7UhLVEWa0yZqqhi7iBAU
puuKTTTJPnOQ4ai69PM00L0Goz4GN0sC7zpwqPGlEv42lvY449Lxfpn1334+RzQ/nCWk836uPmTd
Cx/aSphaPTW4dlZIXPRqd3oT6hll34gE0bj9hSj3NvIVaJzKIQ0s14NnMrwVF1g0x3iiiD4Lo/Ho
fmz+BM51LVJRMSw5Bj1fTrNzg0/r1MossO/b2jAvVmrYisqNKRpuh64tpHuuvWfZ50jDFVDKjn/s
8r2/zB2Ki9wOwmaQejwZzpgLkfRhDynb1sbg5ReBhjopfHlxddIZHxUVweEW7Ptahx8uAiJE8Y6K
qUE2199Kuukw029sRN9ud+dDLUHIp39wz9E6daNzoVN9VyMc7jTy6ZQgS2rzay06TwbcawXst+O6
J7Hwn/BHl1YM5v6MnEUGclp5Bk2PiC1mCtp1QXOztiz0ancTMuesVKXOuNAVVPbVZxVsa2OFbRYB
lRqo9LVixfBi/UQlJiMt/aDn645xJBOjWF2gQu7bVUmSdxUC+nF3mCYBFcTsrxMc6/QZ5rTgrch9
lQ5oZrLdQgZzGw0IRQgbRXJjJlOQhWFA4KzrGjoRaYnPTwW9XtAmw575qGyDOrukUTs6kvcHY8Pi
EzxV9jF8MpzEEvOjAUDwrg9H4nkV6sqjTHHeRcFUCC6tY+UpUExL9aJpI3hs8VKYfQHbyetcDNx9
bxv3IAy3IhZfmfvTEBrzoK11DA5fS0vcJKRDCXqElsjDte0Doup7YagXtWKuLKPQOYgywaT9F1eo
C1WCiuuDwc858r4yb7Fb1TXLBFbR3pXUIxx+nzpKc6DgDowRSUVrU3/6zDYvR1WSJeK/F3pNVCFd
iv9kPBK/aqf5B7rECv9d1nLOiWRKKzeAEFnCGp10Yj/Dj56RfmvtVjU28IBStaqGaEuWfECVWWBx
OvrwEcSXFpnrIhJqNt0S6wrkpY4EBMjdPP/OWbQffn+3QKuLV870g3FMBstXiJ7/pzHpPfCJ9F9+
sbgER83IiIvjpR7ky4C4m7Mt0EJTIokhQ+BTeO/S6/bejZu2QyHe84AVuYoyTwX2lXZdLG/2K7gp
e0RkYcBTc7S6ju1BG9PtX3Rev3FE/qHHnIS6djXFggQlBZOs/UCOD5QtLVOLkmI8cT8Or256ANxS
NSTNkdHYz6HkGrmlhoApqSkxv7FJaWinvZrkNGQcjW9rz/j9DLfzu4GdHoNpfpf/JW8Iy0cBu9Fy
qhWliekE/KnbE1Qy6fTitCtJKBoQvkr0phZj3Pu6nO4B00EaIs5lBTVLZCV70TWtxfUDY2BSWrMF
s+042ypsQgC0mRH4Qoiut3NSegRCzxeoVgikQY2bQO6xSOHl7WXggl2kSZWC7f8HeyB2U0QpRHBQ
5D9XtTwcndLIFtKyYQpOYqo7ZWJNoMrYGK3x2r5Prz2W9HikPqvLdHWfWJ+6y68eYlYEv4PayBxA
jqI2NHXAYlKzX2O0XBdamkistRNYw+pcwL/XkijTNQ+Sv+gHKlSrn5lMyobyMow0kyKjWKGtkx0n
Fp8v1P+wbPDeINlWXsIf66YTHeMY9HBBNiL86TQD96mc2bKk7hBnO3460ymHGf+dGgU2qhtrkTym
R6tGV5zKJGPm5W0POL8irMTOkti2T/QsVctYqByJ0ZgG4kvOgNXqukpzEla9pkRDevKSS7xbLciU
yf/nSD7h0h4vctIH28fHYPO+iYNn7nPcxZp0tLZA+Q90u9ZwYWqmn011d1Wso0nNikqjkTOP+KXd
Re3qtMmj7Pc8s2BGJecmzE00YtvyLf4tVHnPNWJFOdnHnHQ0a489Tu2uGL+BPXz3tdwebuOdV/ZH
QabxIJ3jcu0wAKEbWLRkZdW6xSupIp616B9BocY3YtzIGpEtBzqyDKkU4L0iVtza7Zt+PzJzUDRw
2yIOM7e0Pd+GYp7nog4cWAbJww/6zBPX+flQvlC7cYylQOmq5dIwpPBvcyfyNC/tz7a0fPi4+r+y
wRedgCoc9a2hjwm7337wrnGDLFuWOVl+QICveKn95pBlejtVn065SrXA4w+YmJPiai75P6bAoQ1j
+SPO3qbWWEYkgtxU/uWGiysC3MaVmBmmQL2GJtC8oNBmhRS7w1nKd5XhOeMqCj3CwR+vWjerfUX4
ieTF/XBunnoHvBI5KO19aOWQfuJzZw1IJN1unAERWXr7Elw0TMzfXmnoHG5dMso/bLmQyHmroBQd
5Bsht84sVk+yEqiz4jPZ0MfPNeXdPtUjDEPoBgBMu76yYxispBWeScW7IkIqGeNxkYTWyGEAAyUP
q81rbJQNNygMP+b/m3v0fRM1dzO9TDfxEpCl88fwp0J7O/HaZ+KE5D2WGVh77TJTVKnUWWVjSU5I
bfuucVKrGgPg4rqG3dm8R/P46hV8APkHvdPAv2KevujiDjl+ko0WQioT5z1ir8mjyyMOc2D8CvEJ
MDkjzdP+wi8kpb6JIaqXfmnexaYTmFKZhtP7sCTtUdMOgMRv6Mi3/vWfVNSxqVIKSJ+P6t9e1gqr
UvmleW3VUjQ5gyLVYmXkUSuhazHRhib4nrEGgqGmHXb5G8SN5/1SCbrLfwUQtCYqANH4S4ldLqli
Z/F6md7E43fF7UHCLOcNU51xQvJU5M5YI0rt0bw+Ij1zpc00Nx1/VwJBkdeYo61bIkRecUCozwad
luNbMfSPKI+5OA3Y8KY3HJ/So7t2rVNSg+JIhAqE/5NUNftfofqs74iLqG8BohFpps/0pNNJyLRv
PxFzZpNzaujE4g8FYd+9oNTi+4krcHsw8LY6vRiPY7z+qM9XJ2hVv6HObGB9LbVIn7QrMif3mucW
YJnWeS5nf1SmETreH0qsZ6/+Q6B8n+p184NvviiofCHC3G/0xlsL2aJ7gt+ljU2LkZ6a8BFr1F0Z
y6S9fti/5jN38fgLuhbyjozYJpFSYM+HMDH51MGVUumBI06lSASs+M0FMGMB9kMqXXyC3vzz7PhC
NQxEbV/hsbajlr8ul9brweOYWYh0UnYPDRPfdyF6O/imEqq+IlmM771jZ/lsObxr23reZdq6nTyS
Uhk5qknCLB81dZg4MIbQSMpknTv6ilZ3YGcuZk2sv7BCC2olM+0nRSqpBIdrejAuqf5FTUzgpr+d
IhwWIXTSIKib3vpuOmubxZAirm/Ub+ZemyZJeprdhmw9Rc5q4MqhFFmki8AtZZbiVSINj/9bl5a/
G8JapM8ApqfBP5PmPdDWe2KQxX4qEUcccy9ldfBNQNQ5aJrxW44fgK6i0TMCgQFSSpw9vYtBPv3Q
u8BsT4CrpCS9V6EXHtdBLHWPY6tuHWQPGi7/Up7lqlW5EC5NJ6NdnapLNI9V1OvMdqT6au968A+J
N6QQrXQDzyfuLvOkPJXXbrLusOFZQrKqmLJcD511jc3qLda/JMz/OTq76znGaWb2ORKB6IyUnsX4
JW4Sphhh6Uj7zXZ57C4UcDjFNcGq66OClstsExvbVhqaer1sxxeclwt7mZ0wdxOmrWh6GkU3o+rR
8VifFS9Z8fzUgo5VKXbo1YwUkhG5iBkKKfg0/87YoyWnM+7cyMzRQAS6PZscCZ8dyDjucMTO8F7D
egotASyOYwICrgukkjmeGJuXpNn8SgoLve6glrI09hsr4nWH7f6W3vm8hHVe6Npzujr44qFYuIrg
HaHctpVqryY6q3s1Jv+Jed8xxGC2WtB25i6gp6mi2pDtv6NzqBhyXzleajcvn4xWuUveIRg7i3DF
IFdSe5uL/pOKuH19ObETtP/vZfvV7FbAG4ZkiQc8iVA6mtCbSg2+Y5XBKjMyJiVOAM2BmZGyyDhg
NG3Sj1xENBxXf2MIzmvmUoqxnrIJwlgN0qtXZONWYqppaMqBmJ4NruZ81rv87VyOlSguX+fHZyrV
UhAm2aNSpNZ1HoGF5MXpL5lzUMKMIuWQrMH4rlILX/QD92LEEF1QOM113jefqThN8Agee9Z3Dytk
pjxayo51sZiEEyFVFAeDE486q1ipCdoyPZztsWUb61SfbyXlbpbAUCqMfx4ft7iqEFkN8Nx8X/XS
FaH6re+6eFU58FRA1fBgjXPLpp8ZZTekoW5SKYMtgDEL3ZqurwhS75phbV5bXtest+tJfgC0DYGW
QcLcxI/ZeKK2KJv/35qUqVVolf+nGLP2LaTHhwe620Rmyuu3aXrduVsX9VKwVEMg5xnq2ny4lKJm
rvvdm283ErD9WO3XbISDLiExfxSSvKmwvFG5f2+dPxov8I6x01HAPXrv9eKBTB9SwC50kXslcImu
rWTzS4fPCspqmMX1kpjSm0+zvRFgjhZ2ez4Rs/iv+vMV+aC1oyRi8V70goV3ZreJiNu+uHGSHYfc
+kqcKw0P7wiIonMtjQDM6KSUQatptaPg0hOsZylRohwfw79gjEDPz0X95aWeR/xZ9PsMTCsbsCkH
drKvjwYFEVaEmHphJCfR2Q4dH6Y8jrVY43QWPWbak7BEEiZJ0knkFVjBmzHPS6dabPph3blqNUbj
UIrVCP/p/znr8AUokkgPfLhgA74XU/PByiDtvSLrI23tfivdb5a3WlhXjwDcyJBX1+T4EmxO0yUd
AHJ8yJCTW5fJLFz4P1gBH+1Sne8FJfuhJOP1AudGx9qrzyHIQ2O76fVqMeLnrYnGRo8N0IeWkbt5
IRNoXJmicWhEEG65YW5a36QzoxuNxFHG95O/4W8NLLNg9q1ehWUIxPA4VXrJe7VVvwUecWEkKMY5
4INgtccDfEwCAu0Qfp8N6NwwC09hM2VGtRV3i9hnwv/tWutSVc6YUNzQYvGlcxDtiiO0Qv9euLM4
9xiMqUFVZgqF+9bTKjdXNLbaWmBBeLgq9MNNVkcdzeWX10KYx8QQ8jpDEcrO9upFDF+lxu+XKz/k
KnOq35xYw5Ci1a7NzlBkt2Rhg8zXRlf4eHEqMKCYA2bKV6sCF8a7mnGhhPKCMeO2a+qKCKD8HID7
KuOyEcY0Fj1RHOmuKKLdQRFUbMHr+62es9rBg+uDhetIvdZkwdh0o9ixgh33UXdkXgr5YtWwd1KJ
dVrJumclFBM6f8N/JNybl2/P6Uby1nj/hLRV9d/TrmmmFMF9flUetZLjgY4BoKVG5GfB3UMQcyj4
729RZ567pgOwdTzgBpsr+kZH7IKGDtR+qjCQTn/TMJpQvJRho6OYADH8jDkoiiXf6gwR3pEILluX
dQh82Lb9ODOHa16SbCfk1esiqYx5baJhJWzuX7yRwL8MxGQkJqAxokBL86qlYO21kbgTUNDMBLVB
a8xnPuaOBBLBizbtsWvQpfm3I1+w4ba7F69aHO2ZfwFsye3fzKt4lE+jj9tbr1DLWZlSS6TR2Osp
I0vZSEzp4FTnia7B7wNAutMGD4Xti1vE+lVNasIjo/LrOcj+IW6NFLOqtSpeQiLs8JrjVeKgKA1W
a6GdPK8xvVHsBxA+aWrS8koZZgz4F3HUdbj04mnKdfa2a4ChUxyF+/NaRnAQ885NtQq38vZe2B8Q
WJVac0fMhIumo96MbJLHZ9c9pgwl5XmSMG7F3XQ41U5s3f+S/iouvkfp0D03tD+GONA80s1thlEO
DZ2nRNcioEdhnxok9uLe4Q33BhvMuFcGsraUV4CtbwBJxwt+aEyGzRVEB2MJ4ansmRicj1N/O7MX
+gWbfKzoJ+PkMpDo1f7S+JVh+5Kb1dCwxMEea5kyo0/PFjRmL6isyjnVNh5gKqK0s1R1J7axdKjj
yBEOspNs4BbA7/ZhsCqqs1F1U69V88b8JigD/XA4WpSocDfRezpkCoNhys37BKQ94u40vBECzkFo
LBDS20dhEGCc+I1bopEflgOjW+Z9lk3OvWGjyiL6xWwefpLsNBb8HA5HZpenR+FnRTU54RcX8xxa
R+5MgljVfIFe0mxVZCoNPdBXZVuiUIX07nRouVRvv0F7Mwq7Wfj9MNj5M10+4dTwGdQHEvKbruam
2Dh3E7jaiBWoFDKCsLCJZ+Ud7ltVxsvMYc79sRwGCF6jf7vPUdJprNDtn0THQs4fbqgDKlPgKWdP
6jAnM10UvemsQvvxi4bue0zucrwpi5d47OBXlJ7p7ZQMFpaaGxtGwPyJozAQgnbZr+s3E04S97YB
uAqXJEB+LB0N5z32vHvB5BoDUaKQfJMlTjBJIYyg3WbmP7E5JLP8jdUBwAy+Bg4aSNbjWB0epvR2
hVVv/Z9OWIDnproZ7ca3/eFYcjELRDMqmUtPALsLnSriW4m3PHjVwT+yNBlAXnMsORarmo0Jp3nk
nQEmo8Bs8PU+EuNhB4ELDasv+rKX0M5s1nz9koZlkv7b4iJGk3K0KuRu7WU6HEtQJoeM59j1yB0S
BzuD/nQCwNClwEelVsWOUI+T/+TKmQ7LDu7dBh6b5QJeDEsMmHNtiQLOoa5jEfVHXUR1ceuw4EFr
cW3203gINX4Uz4IheYSFUyN6m0Go0kdwyEtFV3jn23B3tAFsmxzIVoG1XTgfOXuW5gyoq972MqW4
A1q8moFCC/vYd/zmnRx22PaTXPh3lvhIW8iMkiOh+fjjsz08h+GAfAgZWwF9L3eZ7/dbT25Mzydo
5UYmtrXpto6MZzQpwQRAZl8LbOhn5vmybnSU6+qDkIySGuVAxGpoMyjg0QpF2L/xJwXbTlZvq040
ROLWB2pX8Mf7UqTVieB7ipq1B36RecqL+DzXJ6h2K7rbzZlFxT/M0LaqHWirhuQqyH3+g7yAPK43
+Ont99BJyYES1AdUgZuDrb1soAwgJk8G1K4x5+b2MIVWFDZmdgr8Mcj2F1izn7Iaf9TJ6ynuRraL
XIndWfr0DkLLyWtN4uOzn5BoxyjNCt3jDHF6hU6nbvFwg/k7NXOahqBO8+6jTZVgFbXuWeuS0CbB
WP4KESA9wn251fa9yFe1JO9AXqgKF9WtHF5mDoElgoA3BPu115DQ7Ewa1NqvwumE9HB16C5wBFYR
DTErbmJrAMOiBOWzbnwz5zc+kMWrW5HQQiupwBhbro90/Y6a/LdUhOydSmUA769G9NDhfktpT3wT
o67jIIuc+Uvo/zsBIeDJLntYX1beS+Ah11mz8AvqDGMvztpENz2iJ5MyzS+M3APFj7n9ef0u940W
Dv5rzmwDJ+SHHqcY5ihDx/0AjIKnpGGn+QRIgMEC3f55DFpqc45J3W2uZ7XBNUNNpRRbkbd79tBX
13RLrZcjyFbvYQmjGwad5L3Kfrm3MFkB6We6e6UCejd/oxginbn0vuplH9qqIjUe4+Zzak3W6CTi
dYl8SyHy3yy3yx8GXTjuGutq6regF5v38neW4eM5Z2Nm9H77nayo24RbdcVNnPFUSk5VIRN4sWcO
qPTUM+gHf7Z2Eefu3QaAwHPrjlztB4WbXJIpOtjsvxIw19gCKC0ee65fmXZXautuAqEH3BM8zIdr
SNxykm9dCXwMGUVLlqyog1/V1c5hitwORvFGJKv0YzDnke8nuwowzrFHYAB7GD4M+HCz/KfoJhpV
ge8+g8zd52iNvIoEqWQ1CPi7V/DHtcrVDb9C95b/OpCjiIZeJ2WItkHRfHuFlDl4WW6DPKqxW5Eg
EH2PxfRWbmI0zIpr7ZsRfGyWgHAEhmr42HLMRgLMJtkcWxdI598GrBB6dIETKDMrWFbLO4NHVL2A
Dl/G1IFVI0a7VGKbY4sbLhVEXsEDj22ytUN5d+pbAft/o0mK0Qm3Gqg2F5ZLrx35tE4uhCT4rk6R
ODr8Wor4De3viKvWY1GLMqQiL9G5XlNZr8N/fTy1sQxM0IlgepMhx7C1WzoGh+9EjrMq//T1JMOK
HsXrAhnWU4uoTjn9yQzMGhmbKA2p1s0Iz6tnaBimapwVz9kyXCnaWPLyNLULw2Az83tWETIWwU7p
kQ7sc+2gEU6k0aGj7xw/nbYD754Pwb9SLvGnkUQgZ4IGmSUUOlhU6MXsiNdIhlyxw3zqTgkHcuVb
TtxJKU2+HyZGPY4kJsK3QlaZmEwyp8KYc1gp7m/hr1sV1o3KN3sm0GJWAVOwCJYA1oHtZR4UptRy
R7bQuCEAZEq6BqFysex4X5+axtF5qHW69y9fKVON+OCf/FFPX6y9Z37j/VaexyEItJFkFPNu53cN
Ugz2xZ2IaLF+OlvfWz9aKLkomX2v9mt7+UBXQMo9PcFXDyY1sdjNCBIRZiOVKemOqtiJESfPzoxg
zpx1702wDpVYTnRJSJRKqFA1NAg5DE1SwnKhUoH6/aqgZ62u3G1HSouNo/16HnHMLMgzpQlHkXKR
DmGHJug6aLp4BrVMhjkJDLOCRTevc3kXr2akoOOYEi6cieBuL+LmPIb7AXn2yvl618ufsmZ1BJ79
Us7ZILXtb6IKZ/36nkkJbSApCR9fO5oScArZRn8AJgwoivByQtcfAyzH9L2D8wAIRBQ/NDdErejH
+l2bWCesE63t/nNTUHcoEC63TYY9FBhpq9zr1YgBxs/sFKIaGZ+SqyKOOy7/lNh0WqTq2eIeIUYE
v9MYFQdLNWbjYoOGu9316BxX4oThazjztx4tv1FqZhWsft71MPAtPqOQS2YhHmVDyoL+kR92/Apb
lRezjd9g8uPBoCGFYdeO4NmQCMLORKbLjUtLkP97eTzjcF+Deg+w1GJScwLrKFRd+BQItYe6kekM
gXvNf9AudLhANm3Ku6pYKBQdFO+NEZlcCbXELhzOmY4ji7Apglp1jBGflEt7VRT5fEHhtx9XFbrs
ZJn4of0lWHE3+BQxgMeqfzsw/Nvg+4PEYtOdiADf/zAn7VugLFgKFIcXRgnSKBAPH2NM9A/L7p8S
msB8926pwTTjkpBvLXAIXuNIIAP7dYgs2i8uztXlboMF+bKlc0426AuXhLhMpJZZJ/96yeGLrMFN
tdQyqXeKEp2yBUihrHa8SPFYVEuo8575g0v/cTHmDzxUdoHK95OctS70psPjPf4DXLlVSm8e7PKt
LyPdswA+fxWsQkxy8LDk4RQ5K7WY8757729LCEJR60xQYZQ263TfsIvZBGmEMpe2TDvWQSrUQ2X8
ohxXks0T5o4Mqcu1gxopz7iWOWSc7YgpjdfvfguJhaA1BsZXxLk3LoNn0Gi7Gzu5xBpeI+5BBWx1
y/qxA2W9Br3w4+zjIzboKpuGoeHQajv21wuRE+QKxTsrEe8Zn9F1eCZiXKX5ZVI6H+yt1BJjkkit
BRXkxekUny7/LZDyJLtT0HLz0EB2tm72Nw5+oPlBdmEpO9feLVVQLVQ71lrZv34ec043XfY9Qejx
2aL6iM/6GhrE0vdzHBtCu2ZVzg/PfQNW12im/d+rwO7mVh+OnZ5U03Wr9V+/aSSFWFqGneD0ZZfC
rqpxpZ5UM0C2iULCU4SjizbzXoOB7YW0cCsjg6TWo1QITk0c8ZhhHit3jPkSf96+4XLoyCvx4qQA
DXVS0n86B4odXaoxW5dw5PByBkWoShL5yo1s1i4ogmDCnE5f/esdTaLTNoR/i4coa/rGYjMX69Q+
REa+Ol+MfuXgu0vHMI0zi/qNwmsj7D6GhlrX5GpN98krVqSuLBJ7e0skI4Coa+GugJgEO4JX/omT
py9KjY3nrn8YUUfFsscdqEak6AeT0bEjjynjYNTEqmahgdfCPKSA1EPzCrNl+oDbnDUvcVuOmfNt
6AodbFyMZEYaM67DTOD9ONsQLcXp0zHK8OA+EHEAHa5emZ45Sgtld9/rbZgRFAMDb6jku5tLWvNi
DtCxTt2HgbFxX7fCX6e+lj7KFGdhezoSFSC+6DUdmLrF1wE0Se0JUcWfOiq0kePKRdHxWNoxFVJ3
7Swyz6xwq9DQA+U9TjgxilmemzYROmbXdDhM3AFIDN4BdHA+TlfnA464eTVfVH8L/oQvMV4/pooq
O4kkJV+h7IRbJBjApT8aNyfITQ/AhEPb4JXv4lziITor2LnBEY6iHaI6njtmMqXxWcPBH/X+cNW6
dQMIiDrTtYMtef6PiOIWFDhqhYSTzFdDomQMiSXbmSPtvcLqyv9OR/Z4N4JQl6o46k0sGs1ol4XK
tLcT3w5XCxZ1f5fbpz0WB1yBpZYHZpPrt50bMc7oEMZ9aeDWSyQfcKWlEg2z1zQOO6w64TUyajyZ
V2jOe7NDVpk2thXvWcZknQcl/r9qYMYcnyx9iRC1Xstz9On0o1XF/O5U2+AxzjwDmMxm2fJYKJk5
3fjSo+Lvm5eOwbROSkFjh6uMHbLW1xr0dIJdWFJ5KoJ2tYPMFU4MxQHcaHFa5A/jUIx2m6VNycrm
vMV1dOUoVvzde12Em9C84wA33kbUcHywo74YBcAMymZEu33hRXp11G6lFE50Lf+EkyLJGTPESN6d
8lTHjeriyRJ70dIAw9FcBxwcoFXIFNVydjnjaPwLjyivT4rQIu2gVBDpG3TuhEhzyOphe/AEhrB6
R3qFbmZHNYdXb80GeKmFb9s/uUx8lUthw5Ohcp6DTrMmd2UpgOGgJYq8ByjoDl/SP5tUVyi2SVDN
aXoCcTEIyNuYcKNLIn78pWEEkPvtBPmE1PiQ4ZuFEA+UAsnquXjAEACkxzshaqbj5O7L18fc9sdF
se91ZNUueelHe+ApmjVUGN+LGG4rRruL7XMQYR26UmyWcVZZzSEywOzqjpc3OHmPfkNyJtSo9DqQ
Kjf5Dxtph5GtmgHUW8nGV9MGTh/dH0FgxE0n7LI3Dj0h6OVF1Gr1rJCYsnXqaA1EwW/bMvXmCMS+
ig9lydmLAaQeJJz22z92n7mZG6fi8XsT26qrS+qRTIaLRM/1pleKHNdiuU/wEmDRd19FXEOHJVT4
5OyF8MUpk9IJef3STzRBB+pHYnHlpfBMK6Wz6BnOQzlQCpkif27+wP7iMYVAi8qArc/GPcrG/Xoq
esf2YsX/wuzGsFN/kXbe8t9mOC6kF/uLFj8AamWexXZibGArgXye4uV6Mv/0KOt8lj+eMbRh54Vq
NPF+dZYA//wS3xTLcOtqaRmUc9Qu93mkkfLxFjBOztWwh/mS5GV4ORJLuZqCsBjZ9a5eQTi00dZ/
i+HpAzzRJUwYPLLbwUiVw0i7GR5IA4ZKGJeSmUz6Cq6NU98IMsHSZ6S03BDy31D+EuSB3l1cyReK
nOZlWmQJHmACCKoaaP1IY2z37rbo3rI/iAJiD5vzDF33qLmeaAjMtOR1UjJlaZwNR6itLM7KuOeo
/SPC3iiYEY1jgp4TEJgt8CQc0xV2XZDD1an1jFiEp2GZVKO5Z+8tjyC6AwNPGbrrY9EzOVU2auBG
GozjpwMIJCf1adE3eV4QDA0H7195L2w13Mlj1ZDjBIZedC6Mlv9yeCUTyfDNbhU7zyKN4ud3FGim
qM1A/PiuPib+CVKhKWOAyXuH5OSPMG92cPEOfpvMdy9eHrMciJSl11YmYYPHYPAjT+3QL+unyHlH
i97yRropaDPGfzpcm0O3cEDtN9od8d89NhIJcEnBPpTkBClXZre2R9RWCG+jM8T+VpR33/VbvdLv
T1QaqMHzHCeLDjMp38nNygof5WmrqgFd7EkSLOE6DaAQNbyQlIjGWes6JE2TjCwJvj1pPyq+3+Sy
t8wvEdqwjJJ2sFXcBv6N0gfRISEINzcPuAXj4B2Kos8Uidlz3ryTZBbrec98LUpGvDFjT2FDEu4k
fHJECWeHiHJW4tfuxRpoJVCmA2ScFUUnaC1Zb1LYIN7hBxX5pc6jBxOjUXaqDICMAGWEUJNydL6v
QBpGLQEAmWK44DOqLH/Ckn8KLRMtsgyFcfyzYJzB6kPmWeOkW/nD1PPPvZ9AodP/az4oENP8yd2O
npAikJiZnXAeSIglUcl+SfVj86NZgrxGbZcbPloz2Y3GlpVyZ/mTsHcrxZc0cCr9yp4eEN5TRdIS
WtGy93HziGszL3FO2ZF4yJ2s8F7bBh6MOmRdjoqm0mPyThxq6h+9JNyVYgatiu+MLeBa/8SpNagF
t/WJ3/9MdUAuXLO5TAHU+uExzt2xbqRPImmzlHSUKu3R9BX9FqcXp9eAiizSLrOgATTaVqCgD+aF
VAoiRRSWel5aejfdeqJwW9OXl7jXKlile2fM1VEAhzlGIB7aDfBbJ59VhiQ/MF6MNSWwvge6SuUT
3ffAEijQPdyv/RN14iwdqtJQlwmBwKnnlBJKcMCq3unUVQXkw90+qzYkq3DBod2I+LOxsJSzouqT
LyaqcTYe5QKQB/BcZHClfFyfhs87PIlOeLx0wA7CVvFktPwpC4O3r8SThQ6uBWhV00F+o2smxov5
5EaFQ7hzGxwnW/kmHnRrIJBsMgz84mb2iK3nlMjHdJQaKZhNvd/GIMOH83ZTOyJOp+/c2yhRj3ka
AI+IIJ2acHIjpRtEniakc3qlRyDA1X7oIJvRGM7S5GLyB8Asxb1nPSt5dyS1UWpr2+DVZWIBrIiS
vl3lppz7odnhMQDto0Lj/Kpw0aW/kxqHSZsOmASisTKpgQBJ7eWp8I2oEw7g0mLKW8PPfvpnpNzS
3xUxe+c+LaqWS+sKvrq1ykivFmUS6ddizq3l/Vp8kMTaJPfqxfEElAsbUmtXSa8YSrDaYiYl/Xpy
UkdtprsfBg0UQEOnltGpPOVJz18Pt8dvlAE9bhZLyLTnnofXRWJHoxlZ/kLmZYc1bWgwpOsQGwFi
rzZgxcEmDUSMSTqd4eHRIEzFECGw57Kk1IpzqWEHhns8V2Sdl+8wk4rEXvXK9eP0IFqgKoyh9QVC
Ph1QeCvIdgzYtNVmAABhBlsyN0IlR/kLQyUfijoXmQEdozvp2xBymlpWYxMhI3dPryLLwpz4idw7
mM0H05FSGjgkFa2hyYSLmRviO+P+LaEEMFY7A+voJpzGKEZvmIT/PbL1+oygzGKXld/rid2VV7eC
nSrRLbsKu/uL+XtfK1WpST33B9NhxnrED6chxpojBWM4tWG2uA153FafVF1jcaLinZtgVWspW+X2
xidHTVw0j3IJ8v3GT8vQSOGzTWh5hzZR22UnK3lt2skLMuEE895MxH4Ws8MdyoZwrEOI9RiPjwVk
yiRTVIxfzLmNJgM2TZMvwfs1BclaD9YWs+J5UiMSb4gK6yU2oV+SY41VaZgFhjj1kiSWgz2on26f
vR/39RQ52xa6gGzJVnCz3aA7Cwz0nv6p6guwXHamDpskzj/S4rXluzEOaWFWWtC0r2D1456sUOo6
BtLl3oBRkEObZG6krzfLCtyP9FDMZy3IAzDrvOqLyJpbma8oveppiWqDyYa79rXW0D+2U/XKlVsr
KG+Bx+PBtr3zozGe8B0UXw6nIHFQQ0Fh3U70ZiJP7YopLvClZ8PDLm9KPH0WpvNIDMQi0tYTtZ7r
lF6Uw5joZmmpd+84or2N20SOFXC8n1A3E0yO1x7hP+TPIB30l+QBOVOwnil7gnoX88kMwnLQjRCQ
0dv2ATtA8sg5ssoW4e7liWbYDiHy5hU8AQvFbBznXfBCkX3q5/ixdssaspfCGNd6PcNitlmpgpVS
YQnH+CRVTiWb9Rl48Q2wgDwF0O4kBvLVLuzBQDw3quiU3h9wf0eIg21abMO/s4Ghy9WYifDP3+bI
Ml0sywO00ysU7zfQ5G0C0yygdxOoIes4aLsE61DL3l53mZXx0wtKLQcU8+h8MstZIIKjnmlZ7Cvc
0Q6rUAFQ9Ki3D80rCJ9TVR659Pgf5G7WhvZa2dyHGx5jkwluCTZsOvBWm4xjbeAtGdxBnE3Rn7ro
D5YWd+voPbVV3FIkXLsVinNfJq8gTKQ3ZgHGhdmkavQLIjMbBVFP35RNiQTSXuS3glh9UkSmkMn7
8UuZ6pst6SKjGlZWV+yTSaicibE5AMy3IMJ/GU/57uZo0s+DuHHJjKJP/8KQftCWIbKki+9/EB9l
Eo5hp7qJNTlEZbpoTa6C8x/BOtnt/rAuY18sQcWUVwjIgN4HrG8BUVEbUkRfpvmf3yEzCov6TF4C
exc4Ifw1rRSTCki2mdueXYlXIOrjPwLlMOx8QndCZDWmtyVXxvV6A0LZFR+b8MQ0a/EPD5ZeRRUA
J3zLyBrAw/Zw8R3wyUu6GluI31u3R5NEolYjoUlXc2DVyEAt/lJTveAIBd5VTKhHUanNgASMh3aD
nQWpK6qbrbsQ2/9k3ZWcKuFp8NeFThgV1UD4DX+YEFFPMYyHjIiUHh3sFw98Nz4jV4EOso6PseQZ
LIpfZhFWGsUV8odhMQrkNy9sA4IG30O0iATbfExNbGk3F1pt83wGTwXWRfrwEvL5nJ1gTgw6t9Uy
DYBQ/nj4gog84x8LjxgU5Zziog7CMkn5OB7L7wvs2Qm+7tN9/kyv1Sed1hxMswLBx6AJA9LhTOnX
ik2epxkhq4jALR3E3oT+pOOBMePKd32CTuTzP7l3a4V90w53dNcupIwE/Q49BYKbWmsSlwW6jCE8
XCdZSMpSEiaVNmAWhrzQeFrO/tPqaVCQXvGakjgwmHw6AQ1m3IGJHqt9TTT9ULr3q2BkyXdgSpdj
cw466hH+1HmShlP81uq53xN6+Dm4Nx8dftGrxGMik1vCawX+svL+7yazjOIfe6zdQgpqXDFjm9zT
Y56kzhMz4q1MBgBaQ1LJXQTDvu/XAkWsZO0liVHWlkXxNGv5hT8vHn8/iOc8JH4PenvepUUw/XAK
YFGW/RsNGfgwZL2jImeKgauwqf7Wh/L0XD2ElnvF2qAoVfVqKGqtJMrfuBdM9vW3UPdukee9YS9v
8o3zm3rUYOVP8JvynqSBcp8vY0Njkb0xAV2Km9RPHYvg6Liub8yg78eRcMU5LdQH+2m9cqYuAn16
iZJoPvIrs1Xe+P4nXQrBMVeIfSXr6krzptTdig2MFYINhxekBPkPU5xGaMN5efGb2W3Z2C+jIx1A
zjq8I6wZRWW9D841Jh2R9t5j64A00ohtmFpMoxpHYU0dlbQY/prM2zxlrcAB7vbtbfp59fZQOM01
RiurfNkUJVahjUjPLKK7bEmJt3L9GpGSeGHaPrUyFwSMt90eVv/H+SmxIyHVFsG/J22TTGByaWDo
n6kNbHbipFJVhRv3WWIJhMA5G5BYQCxqWOFo10kAgyQ3l81QbqYVvqM1KhGVuisGIx+0P7XI+qKf
9jSj+JG7+UHYUXXk4yZ3mof1MDRKWVuIBXEBe1XLCUCKcyNdn18AiABatvOst26aeZHODQBDhT0S
X+Of4ShARWqy1HfthfMaFfqs6FLB9Hbk/cFpclnSaZgfovnqvQYSdJwRkl8gU0npG9DuxSQeqEa7
yn+yzAx2WLIdKFXJBgX79MD5km1MFSE0TQos9Q43Ho5iqkvruTbAHneSSDa/cYY0fMw+0hMXmHnv
gpLn7dsE6UxfUSFpxk/gIeSt8dIj8UV/ZYwD7A6XfzPeKLKwjLX5DymZqMrp58K/1jvsaPqBosUd
m0dSw//OSRFyuMgWyBQklvF1dYQ0e0Pu2iUT7LEUNlA9rvrVP7Hn5Ky66lqPlhIh/cOif4CeEfzR
CHdaOhiFgjZACkaShBPdLEgVnQiS43CiKnuBxdQZT/c1rFOMselLIpoOf6f91GqHeWyyP4kjX1hz
erEmKQ0ZPrxbj9nkupXFwbeGjW3O6ofz9Jha8LutVR0a6+Nz42UvU9/7CbqzcttK9THQjrno5YCn
xIATrO2pmYjuv8Zb6yJQAU7EaKGeDOzfO6/u1t9L0OGMwjZoXrG8FAi0nAUcxw16oe/Hk9VZCZzd
v3WE5dcOjBjAmoY/wZOYpDCxAR3PTE0/vGyCF2tl2RiB+S3hCw16mrNpTpSFxtfHijDsU+s7qVxS
ttB1AuqNDKlDMhdTO1fnrfdkfmrj+7s3qMhrSWHqqJUNVBrkoqT3gMzIEGqY0J0Zt4CMuLHKfO5h
IaDChyfKazs+yIvA6AWEUpHTvHq8xemcT47fQ41JypPty8Dw/SrKQjg4hepH75xY7qiDnWGY82jb
eiGe2dAKaaX1zDedUOJEavkBYqvgWY2eF1xR7aqpBGCQCEoDBTVt0TaCWB01GcFWgFYeLhJTshwJ
sIo3dj/MsugPfyGRKPLGYk6qCGgH7duQ52ec8GX4ezDeLza5m0aOzIaJ8FiYNwNkSKbmlqsQVROK
qAWuIa97iuFk7ezuZN8q6+mA2azSZDijUqB2x/HgEaVXsnSJUQQ60uaVWpmUx1VrY0v3CCnO5FKH
LOqRLUBYngkaioAt4zVtnY++jLxOMuhEv8ME5sqOeVVKl8zhSQk8U0SkxMztOoaokRZdp9J6wM93
mZwQblpwRZcGPbL/EKDi1dUKw4/oA7NrggEfbXk9z0vD84sHez1CNeAChvP91KlZvEotZU8rsfLe
J8o5kO0shRkLEmSGQ/1Vr1Zd+TnPKkELw6RlQwc0Pb8f8cqLAfPMWIvP2oF374PY0HphHhp9gAKh
JO8Y1Zn9dqv74qRPPz0f0J725YeeVhJ3eXCoIOiXD//uTZ9MdcUcMNyxXHs0YzlZRYpXob6UGE9m
8yQLnr4bAxtzV0m1zmXHySdrBMGVTygARoY8M6gq0zbRc6I3VowC/IGmyK9ik0+dB4l38UJmJ4gU
GPDy0IRmCJgqT/ENWAT6TD6HUlWGzmtS6fJ3uPbf29MBR0Igr433/g55a1s0K5DXIbVyEmtpjPKV
rKtFi8+YRMN1D8/LZAapMvsklfnpHxQ/1jF1g5PkN59G31ocuqy+YZ44YgzG9AMpg3WEYI/U6Wyp
j+zatZnxxxpxnm9VtotBbjtR5ZazJD2DnS9eVt2fnWy67xAhJ3pC4PY0Ps6IDgygAm09PJyqnUnZ
1QS9Tpcq8OR0z12VrvP2jE++fqvW1hombr3OMsxBOzhnn3j+oc1iID1oGC6/oCQJ96rVSUZYZ6GZ
W2jtHF7iSiKsLgTOjoY2hVIlKyuW71Ar5Xlr/KFmYLhVjsDhxrg1ZksgVmk0G4WbdukI6o0koSVx
tQIgWCSeMRNZ4DARpGdNIh6eeFAgWYFgLTXPxbHbmHg/pDtMUNlufu+BGcFb0qibN9i9RDBZuZRX
E6t8S3X9vAAfqV64s8w0j1Nj2dmKy0QM11a6Z2VKI3NnB1R8ZeA3sn426HFISNDoQBZ/Bimc1vCe
aZS9FprJBbjK0VlqlFKICQv1Uhm+ZlX2rH8GgdscamNS6bR9RESxm2foG1HQGg2g5uVmQVyDuwRC
Xhax6e19VXVRb2/NBfe3Xpcqw6s/ipmLIOp3YygRywS9118L0kwknlOolwioni6SfPnHwzdMbB4p
PZBGhHWUr9X+FLMrDb3kqRzrI+SuK+NVihax9UFHN/nzWmz9qYaWRrRM709L/FIh1ly7EhSn0PoJ
5cwh2dr+Z9JYBhMvHtrsFU5QEknJzboEX7+2G9Uv88S40fqZ4G5y0PQN2hGpRDl8ko7PXPUgr12B
WmEcifaPAIwt0E6GjNuuHc20xLq3wzTMUVVdLzK26/tcAX1jwe0ih8zT0noX8LxDiy6Kv9BUBkqa
MxeQwQvGO+PLKTPff0oKBquUYsTN/rI0777lesKFQPzidbOPLWfRJzxjyxNL+J0uohqEykJX7WKy
PHSSy+/TC0N2y6tVrE8mUs6SsQ2l4p0GaoBXsKVe1PXhOb2ltu7tU1RQwZjndgrWYa5qyN1VZlnf
5tUgiNaHYLM/HzSWtvd+m8sakpN8z5UwJPGCVwvSxGYy0tWZ/H/y8cBTL0gWv/zUbBCBWj0sEVAp
+RjeugXM5l4sv0wt9+NqEuEuvUw+wioOWLRDupWjK2rehr6LELF7CAtsraFppEZI/GdbR9tyvmct
bV+ZNC+LJp+avp6qj+8FpSUSVvO8pcA7bwplpbIZh/uL8FBZMj3yRBBbRGa9a/su0UHhXND/hnPj
7hKHWAbLkD6kQ3D5oFD+kVvo3f7nf1C8BBH2CgbyIHzZ91mlH2xG0X0GrDvAwiOl98Y8s3qTcJLp
AfMSHnhYeivOpA4WG9kkYhW3I8WXSqqsEZxP6HmjDpr05FSzt68NIPxq0B3hg+T+gIlrwgKfKUT5
8pK95ZL9VXlZby617bcW4yljJB7+7HXasJr45MsfYtoet2vRHu2SYXm7L740yAGRo4KNwa6dYT+a
9Uz/HPqmky9Ipw1ZdDCM1ipSQl2SIAVlVdDPzarIuTZExyx1/8R1471olM23pHm7kafYwc5J7lNt
ss5fZbIZDsHe5k8+ZyDeNz5/2xdtUc2CSNvOCuImnFPfehA4QDk/nYn/IAHbzccdIK+KP2wZ9AAe
WWHA5yyoKI9LbhT9EHNrXDLCYbpFd15sAVrztswnq9hhYstqeJ9F2Sbp0ptuPX9wvPfs34klde2g
/d2XY8eOrI4NYa+F3lWC6Gb4CPz2TS2bwFn+7b6OBAdyfxwb6owkAVYugM9Tiyi4fnr2uYhlqNgN
vpcCf8apyPA1zJpF4W55iFFZwgnkzncarkCkVFlXuZ8vQd56IRjLf/vB2inu7zSdL3OLqlOwU17v
U7uKbvJAxIjC+EKPec8hKsc6G8ISuxuUndwZ46jDDLRuuZMMvzx21K8DOGjd3LjhjUAUGfcF8gNw
Puynt0Gq+FLL45pK/bFuX7q2mPlug7aAJuGgYou4HBEnDVZh7wQcdZASUMhLJ2zWLj31lgO0fwiT
PpBXmGmLYxNVi0HzzSFxew5Lo1ePn70eBpft6UkTsspLvUMSq+Hsig3gRBXk0yhiUiQyaL6/OgdX
sm1ow4DW0XO20L+nBePkpeULHa4uHpZBaA+VmUdBR7CDGMtg4vVx5Rv52BKnHzPa/4VN80csj2Xw
LMlO/Qwi9trKAPW2Nlj22OxNRmJCOrWzGSxExEuCCFnVLoVTBrxO2r8T1Lhv2nUJci3NC0+7Tvm9
WBTN2HZgyOAY2IDI7iaF0piOqXS9jSuN9gd3JBvOz4mP1j9rmKod1gpNPozr/RvLBS+cvcTy3BYi
XgSNhiTS3ozacl3UDZJ4A+nXldfiiPDIdsVMESXjs1q6KQgiuCCYZLpEUwBeji8aOGJ6O0olGVss
RX3xPj3BJfofbm/IXageSe97QAjmGVXZtrcWbMT4sTn44NRaa8pI0jB1p7VS8UkDNGx7TXIkRF09
hKsKwug/llk2uh4bZbjL8DnpHyPoKOwN1cqYSoLx6HbcsQ3CPpfBT4XZE0nBwzSXarTEQ7EJuJ21
rb1DXMuJemCp8dsLRablL0zxn/rgTE0dRpoaQAFrJd22/30Xm/TzHUc+6gAWS8XKq1W47x7rynzH
EiYpdCMZd9xzrh9Jj1Y6KIjj8UfhsZgukPX18TJ6qb9qyrgWhQtmRctiwdsQFJU86jIG1WcaapvG
FiQHSqLFvGLGuKYWVb+d6txycUxI8LyryK11DaR3h4qnLhKWbLLVQxaWcvH+BHUwchiOVxxQ4NyG
fXxe8gx0QtVhkRR0h3OF/cNumamXmFju9uvlD2Na4lnUHmr0Ut8hkrT5Ai8fjtM5u9cbB1ps9QEy
4Cmp525fi5c7OXhH2a3BorMQ17fxJ5gJna0MCjvTZ8geK0ZU3DnVm7ILRxpY35o85DHxXrmdkGgU
4BOG37oTeRpGzLzhx5rjzSnH38bpCJln/Fm5nWc5mn91GxCC1ZVD51fHtpU+6T/c7LKE8q4GmqaD
2Hm3lE0PV0HXZdThy5VMZBhojBa/8jKA0beZP3/PbgPQNe1e1SCZpMiHcOhXSfZW2SGNF5AFVcpU
fKyuNG0baBB6EmPfjwRSkxI1iLk49h7922l/TjGSYGB/n7PTQcG5V1JsdKRQJej5lrUyuwSohaR9
+q+UuVAoQH8qAV74ebHmDfMphYAExyt7FCLbLSAKLWDyEwWqcqHCPZI/HhIb2YRzIgnio5rHNE07
KGHj1e+8X/WS9Epc3f8S9+ACcZz0TPN2wJzP/KooQafAhXnXuUxJOq/YWok5xTPkXQWdHW0zqWZs
ma4KNvg6W5gZ5gG3UBB1XHkB6jZmgibEk9Y+W1rzE4S50l7MlO9gc7aqPqb0aGRUDIcQrS2y36BE
NEb3RnF3Z+rY3V/UtRuLWxeT4+ZgzTDpH/zDCf3OYaarmBnvjyS9GgcCEQpuMnEj92Qo7/SYl9nV
z/j/dGh1N/MO5jhhXGQQA4P2epezfNqRJQXHIFZXpCFfk1fF2HtbOVfD4v0zZM8i6C4gTMXHfkMz
IZpC7cyk7HHcPSSf0tuK/oLD3X3GoKLU9jL5zJhBwJ8eNnBM647OhP+ncIGM5FYGfXyGhsDCMXXK
0R5X2YEGSG3mihLXNw/jeAfUnYyU5DEfnfnHP3ox4g+4XewhvEiqEMulKX/cFhGyXk0Qx2sFOWYu
U17DpbLf7GsYuHRdjuwCsR9Eue1iP1Br5MgamHxaVKZk+Jh9Ti6hqpK5TETAnWsd/wuxCQNEFdZg
tqRKVO9DAWwIpXJgjYxzVsejpXFLy6bXP7hA9hKg4ZB0D4sPG5Y+cf78lNbcXR8Bn5jBre8mq8F3
8WhPFwUmvXvy3zZl7BILHoOtpPqzrn5m2G5SoM2Z5II0e32n3rX3jsmnE14Zm3FOJh9Mc1Edu8HA
/MyT3uR8mAXqhPkGgrUWN7Rb7Glg1BdHUAoWBSmWcOvTWgLY9mRp23ZUx1Tt44yH+wzdwP0W9byU
tRsEqxYQqGBbH0okwKW5oy/xHAN/LGGDUVrkR+eWPmfJuJVb9uy8UttKefl9qM6FroKKZ7ZC/z9M
migfGwtwBQB1BGnKQ3xJH9KkejVP0ddde5+WnRorTbJyJUouXr0qe+fjT8/G1tIPfG+5ro+9e43/
Np9TaVWClCHq4r9Bmvsupy+hxgdmQ/C00uLVCKF7LtVg4yRzV3YLW4P83NBuX0OF8fEG1gf9AB+3
AZIbFE69+4Uv/HtCrH1xR3OQj+jHBEj/l8V4e52KhwKs7TEFnWgIggvmTlydO9MD5Ys5A5jE2HmC
DN0Bc2P415RUPtthmk8j946DZ/SpaJ7C1LQZoA9RojVbBq7Sb/+3D5gprhxAaT7/kTQcLyVl8Kgv
v/tmzOI1xlvsQHGL+nObzzJarAXDVMYQ4ExzX0zs8oaTOFhnFHBQ7jL9KBOjIxf0LsAADP7bNQb3
uia2U8b3Niw1C7M1t/XgfYMxR6Ko0Gx18AcHwn9bLOhOF9z+vhEDi4M9elpg8pOXu44buQaxda4K
F0jmd7ul6TUkeN2qknSZDxQO97UFh26QM9Unv035Tqoas5Pc2FDapojBWgtq40Rx3+5SH9NKYzUI
RmESsvq3oLlc04hF6tH71MEQlu/MKA+aaEdnPVyhmxrF+9qqhq9lAdDk7Qwa10wlhKCdj0mzUSmT
w4jUdn7BEhzGXCyi6gbQdtGV8cpR6QVVpRFmwnd15K/PQWpB+t2M/utH/gSaiGcolmTE0zawDsYz
ozTPpWpTmoObHRMkgmKx2FBDNBlqcOtxPWPCpp3V8Idxr6T/2WSOms8Lnu+Vc1iX6W6up5CCVnHf
Fl8hZ3FAl75K/4OSxAM9dVp7zAeZSGvQ5ZIPFwltfbc+YucC4FyILlwBMFkn6Po3YkwlbgaHcM75
RyQBVCgnonMBpnvZSAu8xG4xfJaiog/r4x71MZuE31rnh+V3fcbyst26LJfMYaytvZScmwSQ+KJJ
8iafzeaACTPEyGLzAjdnCRtOtApDvbmTceK4cnwrRSxTOgDy6EX8OMAQz/hOrgNHaumPS/ANQo3s
FpQJcPcL/iwZK+fp92JagPPrqHmgVqF0DIU5CVICggWVy/LMVRCdeGUKceWIYmReK5n+YFXxPdlA
QePEGOgXRydcEXqADhe1ISrM18JMRZagz0bTNvnuqowe1fRZkU+N4A1H6y7+a0BMfDeAZOy4ZBOI
7pvZ3CGfDL2JkZ1PbNHF1GJcFhk9soUk73pLsR8tQCcJjZVWz3oYLjWa24ND5/IgPdnQnwMcN+Oy
8xsBorj43eVyA7/7a20A1IqfjfA7h2HOcVIDW7FCUVDMaI62IC0Z+LOb8JCZxFPIirzi1daj+qLx
ooQ2KxfqG3sZaXYQnzedZmG2Hi2wTqwShXhF4T2CDg/ccGUnPyz3ZNbERK6iqFgbZCl5lLdt3sY5
8atOP1HGZwECmaqlaDHsZz9KgyG5k42uCwx3FwKsrTXeIhkuMINF+YITBOKb20ZdtCL2CRFuqOJi
a1/mI9mk1lmMgcnvzGJZOFtA5KPQ0uWp1NsWv20/TYRraRoYvOzGoFxheYblQTRSokteWTSRBgvk
29iI6r2rEoOQTUo70fOmbn+O9lPx2ASHiBLit1CTPbF4Bj6KyFLqTMYESOrBo1TmBzc61eDhBU/K
w29EDJNtiPtyU14fbp4oVpnNxivX8uI3DHINaAsmKhzLbRlssXZNv8VggC/ORKgC4XkzCpPxUn0Y
40FFyGO5eeAjnbVgBEW7TnHB/ZiwiupheTmYVjN4f/MRPZnVlxZ9AF3LpagxRqRRgYOBgCadSO9A
mtq/nDCKUIqTJJhPwlgd3In1vUEmwdU4ON9jH15HBGogelqKTtf9iyWsLFF+691wUU7xPzOmwSl1
2kApmgpki6Mt6FWsfWr3tVNUcciYE/s6Q8xM/vDgzE4T4nprBeKyXXjOaJLIL7WpaaN5cUWSAGw5
qa+BOeBl6cqSpRNEaXd9EIcRGm+gvK7VX27J6p5GeixMZCpq/cpS3g6x54esAIV+bGGFg0CC9dfa
8kNSELGOi/JcP9rHmTo1VvDOkSdLxgP3WEQnv7WKLsoLe12CPhm65GIXhZMvqq2E+MZ3zWK2D0PY
zXJuEZPzQnHw2UFuAtYVz+ymEzg0rCCdqA9CJVTxx9UeK/cSxQ6F59CN4d9aGrlu/ss/177yyoZJ
OkWjxjTGTlN9nQLDhBRCKluA+FKbAleOoLxI6tAJqf8hqo3gzyGy/1TLxMUlnkgTtXEmgXHWoMKX
Yc6UtAAidhQDGSatvMTIOzzh+/9rEiEm6OVEG+Uz/Y3boYJRFTwBhKRvgXMl/RjkX0pRjd03gwuP
msC2nK6qKqXtum6Q1pDr9DQqVGq7SWvvOZeKsZE9V1eWxWjgub0gVGXBrCV6c/8wvDcLz7aOsyFz
vaCn97fk2kxShirGVBN55GzQFVhI/V3ldMdPlropOSKBe8/X9ke9uDDbWtdo6aVCjFc4AKNUX4NO
knfU+0SF8DkkOV/y5v6MeMzG85Mi5IvaYaItwOLNRdOol++aklojegpiDYwlbz+QkEmsz07lQV4x
w7Pgje71MOY4fMlYxJbOM5U5O01LKNvt9pKHznYtj8bD9cwVYfoowfow/o5IVd5BU6BUvCdCMMkE
HsQt1Jyt9gIgAXaVPfPKfWcrtxulbkYyTKXgxbQ+oYtcW11tuYaIbmYCj4tVZp/r/aCX0C97P7vS
lOGgp97CcVWoEBrE9+v4i6+8xibZw+dUViJBw2NGqisYCb/fkGTMxF31ES4dfKRXMToXr/0T/qNz
thmnCWoSg5hsZxNYh8vW07Uw7+AnLcWj8d7HiMv/+1DhwCf6Atp1MJd3pwWctJeG8HG/e1IZrKBQ
dFpM1S/fOHRhC9pm1WB1fyTen4LmVBYQ5RiM7ALgDJNqIkgHtw4MJyQkG+2iwGjj/QJrlC4bD/r/
UooJGIxp2Nij9vIoaCxUK/nGaikoOOI3AY2aB78r4zXYG/USRHZYUhOKE7cDTw+dQ81jW3AvpJIi
Rlmfke+woTyeMTAb6rKX/uFi5XcjBs/WtiLl8NcsW8KbXQpV4boD2VCst2i3Irbm6wY36epfaC+9
uyuwtv8PGMhUpjhSzSm8eKbku/34+b9OLC0krGDaaGTE5nPHe8Ox1n8epIfqo6XAeqveM8YHUpcb
i4LU+11Lfj2l86mXli1MZpN1hVMt2xf+P2me1S63gBaawqkGrz+2/0dCbTI+RVOZf448nLYzcb1B
Ydk6rgMnZUs6l0edqpN9gUFAa0E6ZBBAB+jX2NbgoxcDx2CfgdjXT7/O9BJ3fWeaxfQAKm6XdzXC
mXZcb+/WK5LMxf5WO7uI3gLUgTvqNioZow9ttnaJNDOl5D791QgNJCQ+I0GuBf0K7AKClHxtDuFf
HyGrqETFaClQSkOQ0PvNZaEQcXdfBbGCdkf+VhBwg3b7uq25GIi9WvFvtYInMe0VjU9P2blJtUPH
4TWOzgocpsulI1YfzzJUAPOPeyZ6BpGXJNeRllk2nsqxlIYGTwePbsxa/fH3HIcXHxKHRy2lru7n
0OqEfqxTXPGON1h6hDDSgu8DzkhjSLsvFfxN5T/g8cX25by8g7WhwKd9zqCjtfaiy/Ymee+ivVem
Ss5dgbk1KavdQqUUWxxItsZZKhtguu+jMMUyZX7ivnV7ilWU/3k5SpRiT62KVhtIq1MqCG7CDukT
bVQrGcVFlzo17K5gtmeduHU41jScaWYHxYXxcEmGS5mWFjydOGe4j4Q4hGDCfK2aEJxCsVecSc6D
Ytuijxk0K3U6BJKy/a9OSc+d0HCntGHz4vRGfOkHrwJYvDoTlAwTs6LESKzMtmI5UO4r1cLapQdD
1rTFteqPrzuKkfbGNH3tlYJaN2NhD5Du2nVPsddIQ0Idl5Qj3TnLtBC9fG9cnjS5qxE7EQh1pv4J
Rs8ZeOXupA1PWb4Ffqzx/m9q/s8LI7AGLcDKzBn6mZ0mnHTVR38sVVKDmeRA41q09dJJdjCtUb1P
Sl2K0JbGmljgqdr5ZpPK87ceKcfld7pOsYkeZa9CuPcoFRjVyS6n4Yx3S2lgsFPo+BVoFsyghaq8
sw2m+ysbW1OJ271nRerqDgA9oCz8Wjrk7r80ddK64sKsUkYicGBI3lwScJR1g4SU6fQjXuf5MKvT
7RqE3UfuwOl6IEXvM2SbsraujOy5yL64G8BwVEFOdnEkHmVE72z6ANLq6aK/3kvxedd3ietZG6Y+
c89qckXJ44mWjeLtg/4fO/pwiOMI40KTXSSUaS+wE7w85YOOyySQKEXZYcEIjgZieNOSV1VAhFtR
QL5VpgLL7lmaYqRa2JJV2vJc4XO3LpVU5e0dD1B1kHW9VeFsCKO6D4LhBqPLQ6ffq2iXX8gfFEDF
soAuw1uw52VSI1byT7z9EOx70Ij+YfBEnhHwvyH+x91Q4iecDLtWtgL/kg4l+0G2HMXiBg1XWlje
EXr6C4Tck7maOBWtO7Bkl3AnFoGEGGRO68JYwTsbe0Cyl5GXsnud41qz8gluusI/n9rd0kL/8pi6
g2LVUjypbx3xAbgxxXFRe+bjrFyFuYZ8vWXrqVF+XycCtfKA0CnsWD1azndnLWUN6wy/XwrFceXY
t6gJa3mF/EmKuZlLNrpe1vZXH18kh1KvanEB2orEpiQfTp66K//0mHhJHPixUszpTpL+vDKBkJdJ
dUwRJ13MmB0xHs15FMFKpYp9efebGU9NdxNz03f3Zo2xSP3YrCuXRfTEasMOVTkLu/Kh4BFSONlv
1odw7Yx0omBbNAIHBb8Y4g+qopbFCNhfxo78Amt0k8XIW7dQv/lhbo7w70ChhAaDsvouMKRCAWDE
XaXynFSbDFdik97zKXkJswazZDpLTMQgdNiRVvWrqD3h8KBnG2T1jg7jSuj+7pVlrg3Xz2Scz/AW
6r9qGKVUhPHzcZ/0YGKoTgpsKjHCMsuUnKMe8Klf0OtwmWPIYyWJglTddjwjSzMdh94WkyC9C9ys
Vti0UQaNjx+6C8fjGXrFipXDT1M/RRsP7NmpgKhJ772vZdh4INbZVAwzQEMQcDdFxK5N5NzedvnG
mmKw5a9f7xqVgfZFI2JmdpqYNZO/M4qv8BZ7ZHwnaGgvfiB2/6eMavU2ye3xVRgj7rKqUQTGFqN9
rEBaZQPBjcGdMJw8iPkZW6CnMz0QfWUuUsEjBSy0UJHRwO0hBTLAyf5VKh1n4cRnvn3FTrvEFjsw
gAXVB8Dp4HBEwFjN6rKu5DE3Azji4lNKwmRzOxGrrMK6y5bWq8+XRXp9s2iuD8+qGcEEAyFWgXR6
F7vOdrrnzYHllK1xKP9wtz2+GdoNIw4N6NnUq0O/4RE8O6weANR9nKBKnj7mAH30DLhfxj4ebA+K
Y0kXPnKaKhz1Xw8TmmANqyXgTaCOboV16nGGizzTZdoxhCsxD0qg86amh9kqj+ZtuNAhrtMuHG0O
EQ9uP5r+ratxSEKYSdqe3ZRs4gYzpoVeg3gTFyV1BUfe/UKMCwUglJFnB0t369xLJgu0dCO1ti0F
INsmMa9rGFflpCxTb0q8Gn7x0Z/aqVJ2hFT0UhTFw9SkmTpV4NF+kQ281qzVmiLrdfV8ANzRG6+0
Wv9JL9b2pmlMSa6BWEnBRBHj1fIN0krqd6TdSJKasFqvSK4zJdOzZq/tLEBDgrMxv+aFeqbAxYZO
Ff4+0C+uznasa66cl0GB2dxOootVDStXsUOiaPkkEAZnxXdn6oNr2XgactLtgJavHewwSDXUdwWt
tCv0cHUh1b4FYSJk8ctXUHLZuqBXSOsfTGFcN0HOJZAXiRfAWKdmj55mV9vrA4WUkNOv/2tysPBO
0sWFNYQg7rVwa4I2++FXu6ebEfBpkdMHdDrtAslA40lfS65TpCuHU1O2G+eAJ7cIXpRL5m00SlJg
lV5eJmi3u4cRWhiHtsicrQIrpz2EyGZvmR57hK8MH5zbDKMOLsC/8n7iuoPXAnzRtxYLqi9izdy0
Gy2Pwer18vym8hytrQk+3K5AFIms9yAz4hmLuuxZbgs0USr84gYjG/CrXIR7SPjkfLhLIYKUbAQb
aMuuLKVWB0gFrykQwUktbuQw8Efc14W5L7Lextxkl7cfKDxqswKATv/NHUVpnlBy9jUzLcawlR6z
091pyJJ7aowyQoP29tlKHcfrx4SAhexuSWVcWE3nx1VoEafUyZfHzkLbSZ387Ak2LzfZpsafQQDH
Ja9DQCNikkCXqxVo2A1uc1Q7luaWvaA5Ua7GP5JAIUVDQfLjHQzqhPGHtFEEInM6Ma03aDdZ0IBk
MtSZ9SR9OLDfbQt0HR0q3kyAh70Rxivu+LNAr39i3z6nG2QkoEy+DEU2dS+2Sbhja7UtWYd9hfiX
EHI9GO6KIK5lveZQsPP6000e6oosiZb1w3rm6yfr2F0Mc6VSROGlAiorv2DODaULjqbetD2OD5wn
7VfsG3m7+b+SuH32XX8V0p7UWl9UGT98Eily8Q8xHiAjxlfG5qGCEskUEs6xQJ9mBG1muqkAp9Kb
U7nk3i2iP4uRv8xnng7SXG6/829JTxs+bPHHWle+G2E1eIWmq9pKXKMh6kOBlWW1M0xDv7tKIXMP
8FkFoKYieD9hd99HuUwDG/KCt9eQDDZjh0A2oil2Bv/lJaoBMrrEmZ5ncYZtEvJ9ZH2wuB1qWnpd
+YhVuqJFmk5Gb9Z4ZXlwuGZaEMaZVWTOXu1PbQjKyUwIO3Mj68Fpp1+drMHMQtKwiX0gqR5gcfl8
87X5cFt0dbGTdtlvk1j4usveht7U3QVJr+/UPGBcrhSBhZnzvWgRcZqmtPa9CGmUEd6bdeFWhCQ9
DyN8ZcPKcayArgEBPkOt62Gqoiw+Ye+hzja624k3CARp8QsBxwboyidbfUCAetfbhgi/ZiA6RSMA
ixqBifHp0un2Bao12AUuwOUIfdIprJeblsarKmvocCf9LGsiAucCDU6fW+ntyekhdHvRpFwsC2FR
DYugvaiBq/Sf6ZwePkgzuDL964JF4zF/Wh//xh0oTd6dV1IEM/hyaig6Vcs1wf8ozD2Yd7Tj2Ck3
7yNgqTcOVUOEeL86UkZMeSyFe95K3gGRI+9HLvTt60Rz75Kx77dxHO56TXNbxzhdE9GSQHQOY9Dz
pJkChdULSdZ81yCq2t4L71RI9xZS0KewX4Kx0ZvyKZhIBtxUjVPAydh3nSVlVUXur00uNuzKGNLU
7n4mh2iKl46kEJIUzDIm+cmjgIMpC10IBgv79MwYMRCHta7KA4O0Weq91NJq/qxmzMx8XmZtsvep
cJPsVpcNkoWvJEJklMXvOQv6wFnQ1/m2hJW3IiC9EG1QJJPU9lhTZo8+RvafkXYvw4iV9aeT1LD+
h6RE9OgaECDcgOB/3W3XE8haRhBvZOs4/t63dD8AL7JpHOgqau6jxW1qtWztOkFdJgphzEBapaBq
y1DadQbN6ljaWJnaTtwOVXqixC8H4ALw4Pkan6lWJr0XnW/WZJ7octL4WWlK8zx8Iw9tZpjnqbuT
kzgxInct+FjgsYsf59xf8eH59ZZzTegddrUK/lKSRIIIpMMclM3LKnrP9aLDPioYVfIzbL64JEl3
RXJeaHbX4v0TrUNxFap4OgHrowUumBxt0IGdQnRZkdjN/w8ii3E2WfR6o2mn+Z0d5oEc12oYsatf
vPc1i9CmDcVahGAJcudXWDuqTyBtSYe7NW6wYIhVxId1UJvWeBQG/RNFEB7lGrjcDvolzHa1HWU3
HazTtJ9iB8LYmS7dCvoJQv7pA0lam35NVqSUTfQWAbQeOkfMTH4qin5qA0RaMQJEOx83Ek8u4JGO
1svVWHjU/dwYjnuUVlBY/wnYNosIVk6N3eVLUlBF5/J3zbBV1sKHCWRJQ+ZLNH5a75ZGArX1cDqo
tYxCDjbyY43X+XXsmnL4xS7adljWXzrDRxzBJGagNsEPmWSN1Sn7dKtCB5/85kXxVoD90MpP6sVp
DvOktV3EH+Pv2u50nekRudtqVSr+TGK8qPEeom0/5UOS0eqL049gmGstIeQp8FwlY3kxFvaSPYB2
acEcaTz3C6SgTR68wHC4HazhBelgdy0cuzUxe63WD4nujlHqpAMZZT2RdiG32EjECulJABdDHXnN
p7FNPQ/XfdyLdmZmoxGJzVyIJC2+Bs5BHo1uG1FvsBNqfDb64kjYyJ66wFo9fwvVo5xn2jd6guYI
YU2Z46/aGfUu1GYo3NsEKNchxQWYDIrz9p2RYqESKMZNr2j0XEFFuG0SxHUbIi3uiLCubev+xHzQ
QDdtIuPlsoLhD8KtCJPIaowy5iCj9iCGo2MeRfmNA6/piXbRRc2o/YPb/Cs6hDW2GVpdWSDHTiTt
mST/zKPUyb9wKJ3KCMLR9vktNDDO1dKMf+GfyE6nPGv7ulvgM+36CRivYu2UWcydvX6vbQi4sfOi
dNU6DcvEC8c4RYrJe3xDRBiu1o7oJDvfRN+FqYyBOjwzYcdpPmnpkKhPA12aS/pk2Yfibe5+697r
Y2XRDB9Js26Tn3GrUd0qWo5JAAYEaej3grg3LBRZVFkz4BnLu6/POL56fmusOanEnmsLp9oF/YOa
K4+b+iIMFxpuoNTfmv4wkUc2R6KAcH3DIwYb1PZrOc3AE1mQdFjZUjFsvxTkX/M3GamcwMUMoWCO
4uqWUIAgvpETvPbIgrc5AiGwIVktIpMLRZ1E/KIshqaToOC9s6yKjUgtdjOWm/xRH/J3ykVAduea
V5UvmkeFNK9nPv1h5B8aL2dUb3KwLfsfh82YlAlax+PTbPtsbKoJCvQjyECaqpgSLBXSyi/MLLHv
eFCaUnJu3xrkJeu6WyFa2DR7o2lEb5OwtYhW/+I/LGmqnph5ONcbVnjCTxeY3HlTRZuHlrJ6y+gp
NzoCpHB5AyWcOGl6c8gDM49nVILTuTovEoNT4PJtc8FXBKPTuBqslx/xDEcjqrsTulziy3af0caw
rimVZBoWDRbO018NVsZfQTzkR9jV+RBPrPjOzb3z9GgOMyaOh4G2ZToWJFegvrobadW+/9KSGi5m
Y8nTboq8hRyo3wwIVtBXEUNif3GBXRWw6zj1pfjCgRggjWoC516Xr7Aifiypg7DQdveE1qX6fvLF
b00/IdFv3x+KS7gE5lSnsuMFE0yMOdb+g/hM3aQ6MMEYksHHbnaj621VspFLjbonKw/sUL98eVYs
6ULKiazMbaBUw6ptMWADQywFTmrEaWzO+ddVnhDG0/Xgz8tz2DYTM3GrGxy/kARkFOgH9f9iyz8e
0ew51oiqWX4mRwG411hVgFVCrqBXqJZssMViIoZPdjLkzkg9mh8w+TYwy3zp2QyNOPa9KhRIpsCc
28TPG4gu1lPAbuvpm7gXiVxnINlKX05ieSZaxFKA5n5YFBZ+TnybGrmfhZLuQouurut/qH2oZdFb
/vS6659/byA7cowDvrEg0RPuqiN24aHk9/trxxPVVSBRgToCGFiqUAJ5yRZG/L8nkHHnX9wmlV7e
Ec0EOGnoaT4NztXQiGlxQ2DKZ/WlPj1ggEOEGK6tzGETtZI3nXnnK29owYH+W13KsUYj9ZvApa5K
3t8CVQtzr+vxTYuiUUajHVnFruD83Wh1oNt/3+/ha/AX0rFSYm5pSdk2StpNGV7kl7qckpiYpLpk
MfAihrlvr8REiEO16ftxOw4wEcyB8WEr0r3EyS3TReB8NlBbp4Bjyuuee5c6e2cSzUF5hOhTXWBI
AMJ31H4/3H5Mr0gDNqC1gMrjWGF0L9ugaTzRgs/b22SpDF6r7Y6sgFivKIjikkP+y817ZWjkJc9G
ygRzm9+qg/Mc7unWffP0+EHAIEN30n8omSD6L7R2+x/qmG3Hs6IQm7/mVD+49XrC52FGYtrpJdA9
dc96509E0T4cs2ltthu5r/uIoh9kpVZzhpv2WUz0/U+Gr9L/Afo8ra7lGAlGzGFU5kx5DiCCbfvz
xbw4BVLmvARogXy5TambvFfXLFvpcpLHy7IQydt9YaACJjqtKjXEVePu7hHQoYxTkx6qMxaagzKp
AzkeE5CsYnV9w0H7rCrJW/W7N+rkR5TiVXmpTOkXjhX92tKRvkA6+9SO4FkRPMziL4FVuhN8QBam
dkO/e+TjUDOaGAxNX4wIUneNj2iUV8tL5/GoeDLBBJElAX2V8thtfeBMmhuXDXbqjbr9h06+4rCq
KHYG4EBiW9h/2ZVZJtw2URfjw8cxHBoKBfh/tEGxTiGKrD4hCYYrtm1SDopFqK9J2PILtxWxyHcw
KEFr5Hkip5dApc+i/NJM3Nm+KFx2eN1SHWM4MHKp+dhKZvTHi9ibswIE9ob7KlbyIUfKmAzEkNsA
wkAkJuUnSImCfvWk/NXMKzPJfBn4Je1Kvwqz6N+4I4yy2fHFUhn2VTR49kEd1NogxPDPcayR1ONM
KEkSuYoSyEN4h9jS21h2olTvPHfbi8uoXedjchrZtjNF8oDmdJk1rXov+NeDllKaLHLQ1sLJipmN
3H6iNQr5o7Mj3/5//hVouKATZV45DBwjgf+3vlMZW17pP3O4d1qhrEWx4xzI8htaNpNYPW4rDJb4
I7XnCfTH6kf2dmTEc3+aBB6NrKWM+jKL4p92JNAPi+8Q/p7mxMirnsh2QZqRvUxgHlhBXyeHDE1D
kwvXhc2VQa+j3wX6OzeDyR+T91aS1igz4gs+vFPgIMYGwZ3JXzKxFQPUXrY2vwo2/k26PHOJplJk
SUZ9alLpri+hsXz6nu8xmwrisJbSylkfWa5VJae4UUiQHxX/CEtetQuRQfDwxxeXb8MaGXaU+WwE
fpbwjCSoq3d3McwiDZtsbYYRSZPwUg3tR7mXguHdeidYinvdV0RaqGnP/Z66NHGym8LAClvTWn1j
NALjpID0jtHFg6YHnqrpRX3KgdrHubXhT7+zweE71pKu43iqpnx7qigQ+GHbmMa71bbQecOaBpPQ
dlVsKaaJnsr7r8Ln9ijKNRHOZNdYv9m7EPjxYsN+jGzKcIukzjdXJ/DII05ToOYSFHWjxOlnzbxr
zYUwJ2bHUy7DPKmHnuKRDevfmhCaXP95Cyr3ErNRpU0xlCT/hpzq4wAN2vpbMNLSxRvViEUUdtFP
XHGsh/22qHAR3rnywwQTYR8DejdQmiz03Fc8Co3ZWaqsyIdSrmza99UVWpv2Yt7UaRAMUwzyKtT+
ddgynud05YlX5+GMTicF3XOo6lqAF3/GbC5dJ64mjSTtXuq0UblUgfvz8ddG64doylQDozR/LdG9
Feayu2KWiRVtMrIuAASEThcUHmbosUWDBvZxgitJdzdF+j+WV1SJfa+afxydjQw6588OhrgM36vf
17AxKodqSj0jnSKTuJzrWuEg1raLuJHKMicwYRorTFDZxMgde8/fkDPqzbdgDg11eHX5YfmUwkMs
ofsN/3/pRaemSKqjqOiBCfrTYUrb7W836D0NFIZm6Afz3vUqkRN0zNKmnejWuRZCrPubkylmYlBg
x/o31SrG+JkToEWuCfzfNGQr/+sk3Vrt6fxhBe6MdpIGg5F1QFQtiMR3uhnM/O3C9DI/dLeFaMnm
3xHlxt9x7csX1VHM4Si/+SmOORVu2KGGQjSZrQnOhs7fwzZEDmwMdcpntP22fHP1Yrx4xHw8iK48
pnIlaswS3BLn3xcUIEqdr+NCK/sMfUHTf38mKRAyOe0ia9fGy44oh+hUvD/TL4wt/fAO3pjlHBFz
y0x5qGOJ8Fvrkvn11Rx1NeoA/rvpPFaT9Y+vTwsL0LctNwsRbi1I2VG24bfp1D7GCRT8zc9+d+XO
28thkxvRMoSf40i5sc5bl/G9nXrHAd7ugOAsTXPGh50wMHKBiLA0Ef0wWQ88vwiR/5R6q5gJTz9z
myytg29iqsN/9i3wkrzaKbSKr0T7uxgFUZOrTSzy6bDvHfacUJP4DlIAgjDoEagCJXFmIUrEHSkZ
ZOmm+9/bGpASilUWkimavLvWTO5pG8ySbxab6vJayoYYifXk4cKGkdt65WWAkX3Rg713/FNETcZp
nGdVMKAKQXc1cuuS258jGJEXEd3yqgwnd9cc/PAMzPcmTzW6etuKGaCYqnA9TJUZ6sg4xC3B3oR2
3U7ZCox/DRNwylu65A0u8HQH0VoRM7bbBoOrqSgF3kQ5A2KPSf4E9jDzPdvpFR3M+kgd3TwFq4Dt
HC4TjJ0cl+FL6hDHVOtro6gqDJDTF3fuDSE6DuSr2l0wLaOA/SNU7Dgbn8eFfLrH+ZYLl9e2Vl5H
YQtsWuDp0GUjZfMwlzx3/pKfX2wnjb0HUjFsqk6oLX/weMTI0s3mWw3BHxf7Npj9QEp6vwlUMSS6
GxqUFpDDHLHqmz4oAqB7H4iboOoyQLiZRjQ4MCVSTGfJeHtHFkOEiwt4NzdVHLrtwL3Q03wWdKKK
8cBMf4mEleNs2cP6EAYVxR0Tb2KpLwXx05eamYEonLE+/YQSkWpeKfqytDQ8zD53K6Zbuwo1s9FP
T1IjSL+hZRzIIetawga6FaSZatpQUXxaHYJSUcCgvH7aFcIHR/TDz9coN7vRPQV5hpH1ngRSP5w1
Tk0fMpCvKVriqdapYqTFoPOcbwNfZ79Grag7ov7RhEEjL9hhkMw1/l2cW6PKfpGRGDZdBsE0VHGU
ZR4XW7cYw0eq7JQkORYXr/3hkQcEuOAgtBiy/uqbXWrbCiZvPTGyuM0WtPiNINbqm1GbQBicJiUl
wfdLoNxQ+0ZaTB4BW6LTWhmVGNJS1UrnJ8sJalRy9fFB0pqlBnstLQ6mLRWnVYtAVjvd1+wR2NMw
OveJCS/z+TlSBP15A+43Umieuem0qDIlRziBvq/BrefrBq9D5GoHlxEIf1gTs6aR2Z6A1wlDoD0k
uGIwRx6CUC+B+8baCVvc6TUtHkTrfZaLJkKceuvSav0sJaDptEzEayKGX6ylxg3Yfns9VYWR2Ghm
lFVosQxiDEJ9kuroZaXo+IlJ4VqQtwcOP26HFC7chCNZqr6RtnhR126vaXytesuFTl9maez3xgQa
QOynngKImva6nVitxByYqnYeRayjf2eaOvNzFNflUVXHLQ6caBzcN+785klRiDQs/DWPxsTZSoSj
ITHTjtr2rxAKYHh8bIE7MU4X6B/1iT2WdWHronyzkt01Nf7h2mcoNjaEN0ChizlB/FpnsuAQf99N
ZexyJashJ3hxOHLbsAcfv6MhXLqIHwP20j/yZhu4Hb7QLjRbHlf2bkgkDl5xiouxNWm7+dD59HtU
mC1mn8HfyaV9pcHT9XCl/UZfJSBByJks7T8jhJcR1jH5eC2uMaa3w5kZdK5dvEZN4uXPHC3MIZMZ
ld4XDR6OFPi33dX7PGh5CoSyHW9f6hoVzgmTbJZqz7Noh3phTVdhGyRa3+vwA0XWFmKLofuGR+40
APbur8ThQ0JKUK0DoLdZeydLxPcUt+wu9x9ZGDTOFp5ereAtsq0/P5mi2FPkUDV8dFoNVbAVDvGJ
kda12M3pkZLtmVzg7aRWH6oNSOUe98HORKbx9U53BRcMqJTQS170hJBYvv/XZgVlIIdSTJZ+hPnr
2LNFlYDTVWMe1pw/WRauC2rlKCjZmRvK1aGrhfKTZT51FtEy/ewL7jwD2pfTA+8XrwPNW0rsGwhh
3hGpQkiaQivLmfRpLpFgfjCCrwmOcwtVNa1y2/ybYiHnCh5XroC/xIHWY7cc1u/Q6dxgIYMB90Qf
GpVw6+1Ea/KrsTFjl0tg6Yjr+nwh7Rt48HwqyZuecUpoUSX/y2mOYgVvFuOBkfVM2Qv9XFSFd7l/
mbFqH8R+TviQyGbwipsiDqiOvGUzN28mShKpG+5WPp7fBB525k3Wmn0L1GCl+9H9uVst1UhA01tN
RbS3GJS0gNSqiwflMLSgtxJ/uf0F6C1vsNPPnQbrVoxdHn4AoUW/LHjTisyicKN1h3jlAxbbsy35
hmAPXDHLHbTQ6YD9rfYb9CZ/1Y6lg5VKRf3OWz/g0VMEB7LuGZKHCUgkYp0tR0E6W61AEvVNFAyo
PzPkBzmHchea9coDodon95jSn6eIaRxVGXpXd/RDLvyHGWqs3dmy92Z7znqtMhN0vksj62BTVDrs
Ulc1nCcMt9c4fIxnA/bRK38MXcfK6Q875ldIODzHxiB0F/VDn8ItyiVy4Ny83mmQAwKWU1aXud+h
A8OhLwqyyduMqwBjNNG+IZBx/xLt9Sxny4wWNE1m2/UM0bZsW8XQgLiKqdxdQlOscAxT44FoKYTA
3/OQkaVMosnAzpajgTxp+8Pq1+1zew0o/dKU8A5rEgb0O5RyjfFev9CdI+HrXa3chS7x846YC/zF
YRc0QoLPNRORal079foanf45i5ttFHDRzYAKzFYc19NoGdk/EadYu5TKFANPlKr6UqA3YVvjNGeI
dZsF91p1BSvk1u3bCNKQYjCOFb8KpGcUdG5cjhG95zX0eYIMRpLZpkkz2lyC7GJcVMz21wZyZlm8
scaFVJDEKYga81V+3Gt8efkB5UaswL30SgZd6uFfyRY9kT7wv4QvsPDHABoAC6k8xfPo8FIK6+1u
40bWU4FA7Cso5G1FT50pQnYEndkuEDvFI/GWOOheuWKaDEwKQHTUuX5eDJLEHuwgGoUDqO4yTyr6
0iD3nRkR+MtWM1FsRCUa+/WUYWPLm9xyJZ+I6ho/uEHlwa31teQ2uQUAKxdCzRP/ffSl3hq3/5JX
REsOJs59V3yvtxEdwIbTOhFycaJLQVZ4ZcAYcn789BY8EVzL/UiASwPSn8ErN+vGcLcwwosyLZaa
fnd08GQ7niiW0cjZL2im8jxOCT9Ktv2bRrw0xs2A98ZdDKPSNBSxPU/asw0vX/0VABH/WjZrLt4S
sMJq5jiUAE/2gzsg2K9MkJiInLEb3RIdFi9RrkvwXD5BiNl1EfW+XgkUvl+mEyxy6ZYeqcJjZTSD
A2SydvTibIY8bauKEsE7SEAMjWfc0DPAJagvFEXrAvNlX8d95HPj0en2ukiMjLc1HLNsqYdY1k1n
iQXvQmOZdyR0negKXJ/UMJeMd1MywEXQxTX2THSkr95z2Kv0Lv5HZQ5f0tpz5QTQiUGoiSpDGJFe
7haQaY55jNcLpZfm3WeYuEZQdx7m9gNfH/4bYL9gF+elTdxdG7cqhNmVWZDDrQ3Vx5GS3Ie0uXtK
G3cKTjN/kkdieq3dUFkZtATqRR32tXLc+NEvD7/LWFBTdok3Twqy7YSOCplmZVMxmWbvwqnEUc2k
QeFt0rYGSiIj65DC1/xAT4QY/v5piE2T3zv0Cly/GRfRjnhmX1l+ByjfXX1sZ2mxGqb7qvOZTaMv
PDwjPTpAxol/Xm0gHMK21FV/dtgiUV8urkc7oKZ3zQ3Wr9YXRt6+A44KAUzjeux9I4ch1ayU/86Z
BAm6yyHVLny0HYJRXqY2lu9ybkPwMjOxKYWfeTfQPjtnxxYSBLOBX0NrxbLUzSjON25fRF4U+4K1
I7MwD9y/1ymdU3uHUbTJXl6wV3++TJScYrUv7HKI4NJNsbSQ567mVVGwAH9C9yw6jTjWDu4Tl+3u
1I46AgGbtBcekbwe+AY+fS6CEH7n3HngdytkBbVS1A6WbHLpBBulfbIvBp9ZJ77OmszGHWUDtnvt
J00C1i3G6h0oFWLko1ZLm1h8empmCSyzncNQBprJ1Ton5ZqE1Qis+9iEkkmm1SejIEuUtt2A/YpK
xo7uL7+aCorzu6LF1p4I65uBCSsk0CZSSV2T3inVTwGVAlsA2w2m7qlCYZ/LXwYWEycmVeylR1fL
ENX99LI5SNgewPUcUemljOvEOV5fZUWCpwLH1rH8NFTEeX/hMcTLVDi9yzrkMu0+SwxXU57i2k6T
XbEIm45tbWIhlvLpVxIV213siTUxDixHC/oOXxVk0Rgt4qOQY2cEH9JFt4kIFvPN19nOzl90k1Vc
l44trMOZV4jz8Zo0aiIKdJlu8S2yyxEJKDyoDy6IJ08GF/BCJ4PB7mafj7kU3g4FJ0knE0kKTW4d
PIcpN6Da9GV2eIG9xLVpd4Ja7H794wBZ9x5dHQUF33QhlLg+KEqvBw/f/ZqP876b2cO7tQ61nvNY
zRo0joLA1S/dXAN0mCHNATCTorBVz3+SNr0yOCpHv+CjNJy0qpO4J8Qg/Ou2BNDbMZXeWLO3MdPF
39BGp/YamEyOpZ782LHrm0aefW891kYtG14NJU3i0zMDQA/9PGzTRawUMcM8gMhDn5m8+0cgZ1rM
cHDmcotaFsY/s0kKVW3tWn6A6ZTfDPqJvBmyBqCATfn9NpBsgbAzwxj03K1rL9W9xqMXWGzjlj+Y
8jb+D9qC9jQo/5qyMEQ94J+ecJFpr4tCHX7UQiq0v5aX5sOoP8cKwhYRu7+M4zynk2EBBTBBkCol
dB2CE9zKHC+Yj19UhDj/mVcbtlgwMN4CO42WkOHJlADhSHhrUbhTaPk4522i+9+TaNs3rmd5MuDv
0rVF5fqRmPceBzMhtwEmWSdrLvhdQPqeJPicg7WczwtzbTTqn0Aw8cfjljrSkDpgi4Bsd3g1gKsi
mGwJtfH/PFlCvycLy9W6PfaT/6jzv6j5w87kztrc6qgbz7zgT8UrLHkGtk79nCmAOCunI0cM6jmF
wg46BVgA1UqBWLQKU8joSBFXlI5M7USLPWb+ya6RhGhxGwVcOHCbyhzl9hMOn8V/OO4UMaPn5LiM
WhkaJ1H1vpBOQJr/MXu8+dDY6gUPiV4zphjn8pYb+89YVqA99C+bvw7VSVwggPJrKnbdvoF8qQEQ
ndvUrbFkgYWB+jZ4wZIRWHHA6ImbEqPeEQ5YHBtxnvESdXgg6sjAOjfavbwvUmxHyDtUJ0wIqOwP
FSexC6Dia+CauQ5XyMNmJssN3oNjx8DOjyoFXwwiiCxQlGR9mcOMar9r6TTkPJ8mqcq2H5RrLM9a
SgIRB/bnxAXJlSZ6gQJBCpOFip2WH5lLwm2CeAzfQcowNeGb0kqD7DiE0kI0GRWdltQXVR6nknR6
Ft0aHtlCoSlcAjmnT5pyCdRmn/iERHBX0Ffoq9twkz3+hJ60XldjI9x417hJQX5RTiCXu/8O10TM
PU1K3ls6Y4zjnl0LYpfGovKrF3mxy+7pHR+1wiTkAnY1DxR9NfjPfACVLmAPzaeljMJwI1ZZZg0D
ltYVvfd9auQ8Lyf8wHjyR8iK4Bp2gF41idM3hrDKjTwfQgHT34V2ZvmomEaDcCtYZs6ror8CkDuF
aiQpkaJR6Tw3r+UDhlX206UHunoqXiB2nRtQ0wTseXxApqLCS8UhEQgvUhvEpVgmnAdvzylN3o6h
Hjp2HY+wdDjHdObXsjhe9N0rAIDx162aWyXgRZ/Cp0CLyS3tQ+VEx2kQFg/h8zO0KRUscgjXJTYi
u7xa1+COYJHQBWI//oNIfQzvoGKAsAEoWDWZ99l+Teb/6Yu2QH0zACb/21iD0N+okYsYmPG891Sl
hFkcbMKbPfa6INYY0VwsEH7UlD5uWKVVM0gDbs5w25abiqxnQFmYDbwyVTuLFVu6HjDNhBn6qLM+
+Qa9SpFKtXRFVujBRZeTOmNvRphCbcsqNAr0u2fR6JuwbGN4fY2pOnxgK9iaQO63AKTvY4UgaNzL
MokbNNKuvmlxgTNVT4pSOyXYFcLVFNCsF2iNFF/02KJ+WbBp7FFg0bztEtzW2FSoUeN6A1pOLTWd
JPXpAyBl+FNepTTdfZT8+vf+opF+Ps3JHhJ1Z6ivazA+qNug6GKhdTNvIicHzl4gV6sgSulWQHMq
0fwIFb3JK3DX86pgtiH1vzhltuP9G/2BLGuZCX+SWnICavRgcUnTxAxbkzc73TgUJ7M84RBCL+jq
zzXm4W8UnLZHXVzYyKpXUcD3d5/jxax0vO1te08X0cbp2JeISMhDJ0F4moOhYXcyV+ItIbntgPeD
igmA1B72fKezjVGM4ccc9+Icm623vq+rKFKqksH2YJcEE8u443AT2gHN4ki6R3RgLLGk/TpB1Syj
vPozN0ZMpDW096vanfGz2UIB3L8kubWnYs4SNWbRA42DExGOFaZE0UxzZaksrHtKtHvzebaYaoq5
Xqkx/tIXsjKB/SfuJURiK0XE6RYAvbi2OE9dgMDKBq5BvcZjcJBAZQu3QQrMglBGWwdM61A1D3eh
cdW788RaIFuyf02d5KKDHDeK84S89lITeysSSZ2BeNoIr7wXteh8g5AiDqOJZH8FojljByy9T/Nd
rM3UtbDP2GdWbOpUUk42CWkml0cM+CGJ7EvBW/dB9g+NeT7tiigojm5/1FxPgB0svWcCJ2GNcLv1
roba+4Y1LmRiHZZDzOrhxduP/I4ZEDD/6LXq2PmGaq8WBJD6YC8u5aFbxo6uywaUwg7DmXgfX1fW
We2tyYNNznL7ZOVMGf698zww+sxXRvf9RDCZZBXc2wZwkcreNvaNFNCawdk2TO6YgjXjMl3+L2dl
afo5/buhw14lG+t566vmBkZ+1mcVUQuAMElsPL3GrZvUhCIe21GF35ej0sKCr/rKvinToI16ECx9
qFZM8eEYlFZbqGYq/SM0u0xOSqNgKN/2Mqi3p4VsKWpkXkEgUAXkhH+YWQT/CtWW8egtbmJx0wW0
h8OeC4nDdYtjks0SFQkfJFckuuj0Rcs79Pw57BVMuVsZKg0Ov2d87FwqlduNyz452HItprh+FnDD
61qONX51QXHVACnwCFXOwnnR1pJGdIM1h3wEsrzjH5TmtTd+1gn600Gn7Xf0zC6QlQ+DnBHHQKDR
s4HOyMRJ3Gn+3i3PUp2W5bcj+gRoFU+VvjaI2hoXuBn1Cz/BTqBI/Wdt+o4+b6OZ65mWjTyCUmXl
teDTjxQK4egBt3YsnE7lHRKHCdq0ik+EZ2jmIaGGYLOpigcsdl7+TC55LBQATqmXPGFpQpZIk/80
iZV1GCCL7LyKDXI10pD/H258Ew+zysRSGTQRIryt3f3H7t0Kalm4I4ube4WqIjZpxZYxvMgtLeg7
Qfmb8CnU4xRy62WBwRL/hriGqa9BP3KXVRkZeQgb4m01V5V+BkquFePusJv0X2T/sA+KdYNcc4R1
RBYwJSByXaIt5JnF+IXEsfvVCLXpNWkXwVcuFHklcbX92tgSbkoZg5GZte0v85GXwN3ajszUhg+x
JMmmqaAeJ/yGEIqE3a9IaYWxLN0F61JH5wNtwgV3E/QWkFrvrRyBrH5VK3RnGfS1p1KW45WXgLXj
m4Vp6FUbXb7T3TJ6Qh9eAEajuYqpXLa/VEFLVLQ1zMb3FzfY+r2ujQ1QN1Ctu79LYEbNWSn2GJMZ
O/EtpAmKYsXwO57M2EFud7Ze4fhGj+By1kqUpu5bb21cgdHesqOlBNShSAvxjqaSLWNSaJ5O2+ih
eQfXD7nA3XgFeD3mLBoKUGeg9v8K7SjXojpWGUeUQYY4EXTFVz2qUTFL5HqViTsR1lba1jXPWa3a
b/J5Pw3t8plbUj0C9vf/aiOKmBYJB2c/Rww6Xp64OJ47PGKDRhMOkikQw0OfFh4cwVmzWhvWF8JR
XNHRcOyi/j1J6q/YpTBUTKq42Vn6NvtnDGfilyXWl1kGft9hG12YRaoXTy4zAes4QuLNa0vh5Qnq
MCUbGRW7YvLmXXOPLmZyvMSpbsXZlU5FX1AdSjhoaTqisrDAcEqvaXWGP7T1jgbMD446ZiWq/K6E
q05Yb24Ygo+s9rPoIcwbHM6b2PPxQAiv87VGox6DbsTUtWqMkPo+tHVjvoHMVYhLqVCQ2pVCeDK8
D7DYw3cxq+pt/am2Nc3ztU4Zfk6b9yxdf+5oc4f2dZhCwW2FdYF8dk/tLK49EUlWRdj/uPGE+jpF
Y/Ok4W2ECjhxHWMYTCXeLN9ryLuqtpYqEGxZS4UHgfAWKz2M6Teag2hErqMHszeGifVKihMI3ati
Q5LcjGYBnKA6t9Eea5HfDghM6nAAJfV4F3Sspt+EedyhdbIv6blWsuqQcsBZZ5DYGp2gZeeEa/J/
0GDz/l04qpRbPW7wn+j1YldAhZsgtYoK6YP31QH+w57EKPyqAbvKfmRUzbbsQb1isvk7kuy6L4fE
pTq1nwweGGtelXmKiSJp7H3vrkOJ07sOe1DCxn0Z5tAneoWwtGyRMSy2djjU7uNWHIvCRqbTeQRV
HleK0dlwUp/5xDYO2/JMC/+iFeelkJQEUeHVq2280XvvIkkN4WtpFBoJDI7NWo2YOVmmkDbkvYmr
TYGBa5Pzi0qERmicBeLkaOQYthZqxNRlbkvgUvTEZDZs+WLzFS/fL2gYeTQHs3AKmLrXyavuhfBN
tnkLnQpZMEqNknua4qVal0nvKc6ssVXoBjmGppvIR3NNWD7pg5WzxZ7aJRCynGLEyrnvelJSq903
viKlSq+2rQchMZ4R+e2ifRFN30q/sLLXjHz2pae3zkCUhHAAFMpuroFJgQIguCVfWDIFTvUpmsPO
RACUN1MP5zcTksHu9cnYknzv8bK3Fxkvr2ztygl1J2lqo0/l1EJ+Y2H6I5TUS85Z4D4qojf+tx/A
mHZnh3cXcGe2B3tK2lEQMU2wRmI4YvsrqvPNSTsK6l2fDUiF26ZUNxG2OEtFNKARX3NZwP4EYqQ0
r9TNPPWlxkw/jByPNn2XB3fx95C+67o4SkPMzMO103lkFpN0dgBVCV5gTBVC+TJKtPjFUCqoj0v2
4xov56FNWrSVu2Evu5IaRFa3Rc84nBLmxh8PVJ2DBWeUM8DygpERLHDOgGJi9gY/HWWibzqalAzr
37BfN+btpgtyaBePCZlirpRATft2/C0Kz6PXmlrVHYG+Pe/D1IntIpeSnSEEORR4HHrKy1SziS6f
fzx8QlrvFsgGl06TorViXkltehx7lwW3rV7t4zzAGQW42kTX2OnvLa9jdAVYR0jXnMGD9cmE77gO
sOdlCKgg9+XVSvK/iCHy5VEbXEdTaWECnVPQDCr6gGwXHLCxvoHo7FXbDxcVPtCWW+FQQJU6Mbui
IEj34nMcX5cq25QDdzGbPG8+bflT6An6bKy10dM3IAm6ALF2WS4j2IDVcJNRO9c1baZIBQE7+h7x
X5hJvRMoeAIJSuc78Ss1j1aj/BeU3Yh0i5VJHQ8nUGqebQDQNGZ5F/PNL6hT5JPPdnUYLt4K2dx+
6Fzcgsc368oVV5YGbOL+1umJDSfreT1GZpA0iMzmOqGOJdVgDoe+/G3gC5roYHoiBjfFCmnu8Qn/
dJ0GckTRDaXxdkTwjSto5To8YAi/5iINs4/xF69DyxYjEOXnQZVW9xU3agqXBKLaAnwwZrh9xbjD
qZ/UKmQYDODWRyfPtzymi2rNy7KGdeh1vxjwnHIrxbq/G6vkw1DYRin3anq88BQR7jTG5t47ApcE
nGhfSxYB2utPedSNxLnFTLzkP7/KFrEAuUDYvzOgmvnl+q3z5zB5k8m13l86a7PDcQ3OJqJEkZSh
iWB/bjQ43pZIm+jyzhXXgi4U3d9JpG1HGUvowGzMjZXSbPnXUiO59zgN83QCiEwiVnkcFzC4fG4E
WR8vVEJkqhFLa7OrgKNrRF560av4Re2d597khFqnvN+3EK6Qwtw1q9r4KsqZuzgU8eXsJZ/tON2a
pnyEsB8zx2nnAgFvoDghjKD+EDdqFlC8xyhQDgk8IQ7Q7iy5OQKti+HwuXhMeM9CQ6tAQ4HclCRZ
mTwxp6zjb/30efN3KJWIVaM/YwprOu64mbfu/bzzib5bsXBc38jMt5cx04JH76Lygy8bpXI+d3J2
TFlM7szjEre2JfP9twA8lIJLxPjU/jVEak+6Hcq4H86l0jX1+rH+ua7rGNSvl4mqvCihhCHikAWv
RGdhvnvx2bngajHyevmCXO9Gs8mXMTHuVtGCktYS7TMwqEjBNtraKbvt/vC8R4ZlwvgQu0V3VHcv
8Q7/FOwkert10vLjyqSDvcLTgOu3k1TN3lNwYL1p+ICY8eQ9kfCac70UuMVFE7tFisldZK88llXl
Mx2Jdr1CGLlOgQ1EFhbMoTa4J2IoVtOmK7YPFSgc3UmDix82pgkXa8eZCT5m2QUN5BAAk9+gBCir
5u8TDhUpGKIJWcwYZO+Z3PWF9cFj/iP4kfmf642yN+6UATpe712yb/q25J4a4+Sv0rUE90nUyB5C
QuMb0wNIwzkQzw7Dcmcf08voRHeRc5cS640pD4+E9X+UIo3e2B/X2PrdNzw8lvkm8eZUD1txqeNu
Rzymq6NChrq8djEPzQealqMoO9ixpuQe3AvoUv7MDmwOMdrkxWOc8Xd+aNRx/pth4Jc+z30O96IG
13x1RPzuEjHmB2k/RrLuF+mNLIJ4d1H/IEqZoSUdtQZlm530Zv1o58PLyn9lhGQ3rHUM5ScCEZaU
omrzg4iqK/H+DWoqFEptzggLPX4ehOFSV5h/2h1qf6Cds3l+IZ3U+9BDkbx6LTFbELWtoQ05ea+R
EO+XaIuqkf6M4gVx8sZEG88UADa7K0OFsMcBGmv0shCUJsiSrZIa8yRv8Jvcue9Cuqyw0lFL85Ok
KiGenTmIzOiJ82g1sGkf2/Vu5WnZuj5IzWVXUyp7vRSAuM+gizW+k/zvln+QT2xBmvcwnNKlzUhf
5tCYf333jC5mB0mP+EdA1CsQEAidXkvZNyVPptraXk/70iWAtAeGzLoLo5EH+QCgCjv7EBySd/dj
u7lR0IHH5pP80gOt5NB/129NfoobzMq7Vm4rh/cpdvD5HJU3c8C9+PEgtsCfo1r3XtjWZkI+oymm
0bhvy0HipiTQvuriGZikP0HcjovKyUDCYpXMMJtWoNZJRAJ69k0X0AbE/V8cBHWrecvPIrkTU/Jz
WsUd0IC3l6uJ+HQM7DcW0qbDe2jCcSwIsbkEjPZRv1DY0NWtC1guW4t8wUynzOI412uoJyDz/E9H
XgxJCuUACm9QDJV5m3moOIzJr/VrCGQ11RMwdQS/AdgF+v/h8lmuCGn1dw9FXsk7cURfSSzZSei0
CuTX9O6QSVrxs8uWrUIdiV2WCClnYI5ljcX4eNK8FA3o8SKRz5aT54znmCRp9TIaDRYZEfhCZ5Gu
Ev+v9gHLcEl11fBQwgGUR9kpD2VBfF0BYJVCsXN9DPXz3TJg9pSTwNL4m7khENbjjzJ7GAebaUDQ
Yp1ZSCz1Qrjcrn2gxfiLkSnI/olBURq4XIOe20w4Y+cpcYdqmsQjAntf62LSMTyxbLI1qVcMt7eQ
T10QuyX2KBtfwOAgGDcZ8k011LugqVQQV+msS7s0pSIZWdMoSNpJuX3J8cymkusEDtFzwrqt6uwE
j5C4PUv2oqMQKjIggngrVa0t1qAmrIZehQHHbbit/cfehm0IOVUVkxaSYoAitLCR34Hfp/FAiVfk
/iGylfZUlvQDXBOtaa4LXiZLJkpPLEO1qd4jEQvRV95bGjNnxAlI6ZpUYcJJKNlNfnUTxnlIYSYj
TVaDIoAUkH4EkEfPJGGiINpq4UnnrOhWbKvO+/rEmq240MLpBdTCA/hhZCG73Ce31D+ZaDJPnGpO
jGqmVftzia5LyQ2RjrLHSE2IwLn0Id+ON2P8bpp8AX60opBQ0RVbuMcZmZrDdQJyLjCf57H/OdXX
jPpgO5h8n4WPZpNqUfwfqWPMYGD0izZypXs/zL2BXijpEeC7zHTxiCU4wWMgGTQFpskbXECOgK7C
i9cG9umPqMQ18JGCN3IKH7cqGRUWtxX033fRMcAHHrcLnQobetpVENRooCr9v50yr0ya53NQfrUs
xAaSa6gyDfJSQaUAQ5EQ7IeSRL5ICHI1c8u+fET+LhhpiiWLEtId2sINcjhs2CrJPx4qnEDY7PmQ
x8/oThIECAV1qilJmFpCO70pp/IHMMyxCPxu701qKyhEa529nR/9CMn2KZ8nzqC0/PXsAmQKm42f
gJ3bw9jXrXNmn4VWGqLaBox+BvZoEFGRhsnRAsSoa+/BVNPqEwJTwX5mMto0W/hdZUGj6IpPkR6r
eQ9Se70P67FuVmZSTAWdnALyxgtcnhvN38M1FRjk0U7vYCuehT5+A7daWYBeen6gyjXpzLuyZxib
Womc0wKty4UNy15t2xeVhRG2WKojB/x6iTY6vj6Wg31HbXgp93eZm51xt574TDnuCBQtFtCNXYn0
n/i3BplIkvkoGINKXrXDoX/71+jY05ZjLWSKHj9CnqO4UUDqo83NKOoSWFLTVHXUCyAy2phXOhLc
Jqn7odCt/KmjPoEU0BGDoKaxjf4aHmBUgv+3Q+nZCm0FNcabA2skxuNeBxAnPSPabIPgJyyXXSrj
AgymySxT3hpaqdIdML9ZDMAsYVIUJdsNHFQWqSqK2E0dbMyszV/GbDpTLJ3mCcdD09DygOn1wXOj
hWkWdU+yluvyEMAlnW/4n7Z5MPMW7EI+hZ5mOJsi+zLblQtJ2xzn7x5u6+jH/gc5K1+BY5D+93ur
Tl9GHjomYZnCc5hn9sYyBOQGtE2sj5GHq5Q0/V/hVM0s11j4ZlmXjrCUU9NuZg3iftSLPrssegE/
GX/0/XaWwaZS37LHlh+3C57IDuL7FvIJp7JZdjrkHx2M/U6wxAq2ejCNH24h3Xh4TU5+4Fo6aC1e
vMTLDZAK8hpDVbwF5XJ7jXuDFhBNzFXnb0JHoox630YIcc8x+SpacjTwtmiSkYbhefpJ5dDnZXqf
dZI7IcWgAqfbcLojH8vM1e/qWEHeNADFS4b7+C7S52hyy19HCDtXpzI/+7gWJtiDZrQE6zO6+2wY
8bIKcj1+LVZQxhDFIC/LgCl5vFWrRxDGUUGr5bvZmlH1ECdLEabuaJnxI3hUv/6q8GjXOB4LvXhb
pYYe/dPFMSH9zHa6feZY0MT3jntQiRXVj6hc5wwvg4L+2DQoAC8iSbXwq+RevQ1Pa9W984GxZxM/
Mz2X6v1KQFXHB9HFy+O494eIXuQ4xhKuwVqEMybpGnML68ZlZR+MZ9pwkG8IU1jDnLWIKh8/pj9J
pcY0iAxjx5Kx9ilJw7jTT1hXKg9dsGWiWjM81gAnQ5OpOpGrjRq/oQtzMZP+kwufOgyogwfAnFP3
NSKw0ZdbE++xwu2cCr8BAphYnS3tXpj66xR9AVns7GnA8T/mG9XRgwHTPQMRVr2pgeJKjI6SKnXz
CUVKs7h9ZcCKp7LfjMNaQE/d7zkkEqfOvTBPeFmuLdQxKFzJndsMC4qebLy4yVPLl4YfGJWvACa7
N9pe/up9wW74Ecw1GwWla+0kZJdLbawEYc6/mHAuWpFPozaYcDIws3FiuC8rad/GBhF0Xa0iwckM
I13wMHg2lCzV3L8F+FgInNzHDoK6faXpQYtHKQjT1QaqR0vObP/dX1JQZXEcIamJrpQIWs9Wb5u/
x8B6r5FBtkgdTi9X5nv8iHC9OUQ2vTKNYxVz6yYKrsUyJdrd0OE3i1o3MqI5eA89pvWfMyGFenqX
viCxiqiN9t3eDdr6YKXfxKP5ig46wlQiyNiFt6SS2EsSVyuOU9RH7ZbNAzLMlauLq18Zy5eNLZcB
in2ifiI+79OGD8dhfwwRAOABaXkJl8cW46CEWBZVYZkPsuSl55LZJic2Nl8AvI6IkUpcYhAErxrw
ygKGbs9dai/3/GzkOQ1o8euNg+/9twWaDKhdf83xKTX4bFJbgoUj7TbCLfMSA4MH97zcF1wf/HbJ
nxbRMrGpzuufiZu1UnksA8+VXsP3lhFMQJy8xr5d4GLX5i421VgibhZOVYeH52vc9viLiwIWuQIb
3krJ6lYg/n0bJOym7uyqJ0b+B4nx7PlRUE22UpOYGIAdgsJ0nEBXtla0SdUTsZXuufPLUwFcThC0
/nV0YNwmFRw4u+t+HgNqfCC+XmHWdh4+KYeFBeOP8Yer2/lhEIkMIIhii+BdhVZfEE3mgeKKWIHf
PS8iRTipCPSc4T7Bk3XXi+5oaVd6otTnf6gZQnitKTPbdTivWvRFMpYlmmqhgJqvhLQFsGL4fed/
wLsY+eCS3H8+YK01ZPd6nuxrB/yMt++k6hCwGLoXtn5d76qZlH4/6ZgdZWn3GqvYaWCK3fJRfYy1
RTDeN9XxyaFJtituoMHdfQo1BYY2DRjXoOcmeWfp68YRkANDB+OOgxGX5ox9SlGZFB69Uon1/C2K
N5WtgMArcE1Rcv3KFjYRRdZ/I+kSMi/+83sLNowvjoXBcuMuYNfj3vyKrSEIzwF4C7GoyxQzfon0
+xiTxwk2LYnM7aYtelJirpkGpvx4eYSQtu7YyK4u7D9rEhmNDEZMabkH1z2gQJj9cymYmt+xj6Gc
mnX8H3sdUzWX5KzkSA9Tsh5wbmr73k0czZ5tfTtoG30uBd2MKvfEocc95KyiRxO1ZR9qDxepFE8r
EEj3JGYbySASPglwBz1YaeMGTGtlRmHnMgk6bh98oSo2y9UZZfMcQb4Xy0QKBSIUv8V1L7z7Rx3K
ZY7pPM6yIvRE0BBR+I3cimF5m+JtvKmts6qWyust+PeWyJB6+pZtpmnAx6yNDg0jjZ19i5RtdFDZ
ORzwMSPNzl9KSU1K+t9+XJ/yaVWNLjGbj3Xaimh9/c7goeXhzWnzOiNOus3NXOKf3hbBKtrYc9M5
uuT3BmEZKrHUZKLmLO53le+0StH4iGlyNTxnvSWhAw0O5Lo4qbmzZ8Hj2L82iwX0SGjoL0eK741f
yi0hEnpz/286F95s9MTy41Lrlc3bGA6Af6bbwMyjwjppNcxpNxH9VWjwtPbQc5W7Wn/f2Rh2V/P2
HdfYCG0s2oOxFm5hmeBdm2/ttaVh6Qba0Ei/6ayI/lxnLY1PCIFvRX65BcycF3FqOhOnTDKbrOpf
K28ab1QrrWAYbUzEK++H+qwrprxnQ24+x4ObBEgeS4zAmsJ+Znlkt6PNHBp/Pzntor4P8/tYZAG8
cZP5iEhBJCa1YF+134mXVon/JLLW3aSwcMS9jj/PK+nKlvfDr47LXmMxbR/4usED7wMTRz1gRcf+
caE3tvl/4UYafnm12BD7t+vUUfJQ8vSwdnGP/VY9ugqdr/p+VFLDIStM4IcKNmBn8CFSsS5DB/+p
24Ur38LljO70Wi/T1AGQdWwV4sIak0OvBe1XxekHt1KwSyIxzvTp6DvkzjvEhPw71c4/om8nbEge
M7YCiqLFiRIolYKXTpnrOpeikr5oLzS3AcHbIwx5bFjVk4JHEs8HX06EykcHnuj+UNcXOo/NJO3I
p5sE2gCVC+ZyM7+FhnGn3TgtArFq0I5FyxOqEohmebXKpyXTbb7WdnqpxjFvuV5eQgmKCgaLK+5x
qHbPvuJ7BSVHAIkFPZgqn0Qdsd6Qqf/odFIxXi33X31cT3g+d8tCJ6z5tUuvJJhD0ZA85oeJuk0f
5jg8crNGG3si3W8x2xgcV5ZVjipST8ATSwL49eQdDeVprjSuhUobv256hFTsDJOJwtVDDhuV/oyU
CJMjk08sUirJJWORcWNBz/iNep9vCCqXbrC9p8f+8lUW7iPlqxzxN1B7SM5pWvyk/M08I5fmvxs9
3pGcfobernvHwkdoQiHFr6edhh5v5VZygHfu3sLaKz/qjq9sId+Y5m+J7Zz+9a5dyVNF9RDJb0ib
viwt8erOZHNXSX3sr2teCR+tOUA1CG2xp/nBlcsAOTWPJfKmvuPD0112jMXv6deWXAuGidzZUZ0S
KAPjyRJJ0ffsddsdvmmGKTLRWbppzjG97lsbBOgDlnMY4UCqVWurlQ0mMWzJ7Bm1/QQRwk1+h26A
JK7OgOarlQMhHRjEcMr5a3voJ6ZwjCSaBYrB9aDzhDZV+hjrjsZrbmmLlHsHoKTF+p3d2d6F+CSB
X5eCbI0wQhRno4aBmIfd2VnQFwHKWaAR8Rrv3bbeUpz+RHs1/9Ibw+Y9VQcrk8EppgnrMivjsO7V
jWRaWh8pJ4siem0z2U1IyV66G4wuw5OOB75Czx4VvHIn7U3ns7KbMF7hAA6VCc5itMLl2TONLMjz
o8hQFeabz4IBBVruP21ByLZnpofF7iNdrLW1WrTZILdWuujbTPQna68lg2KQI3+0GnFejC0j9zWv
V3Q9q/p1rpppztWWrvCu/bA1br9LQfJ3MofcJUjek5q9Eg5NlGogwFkHxR3wBcIl/Xm9KojyNPrs
gMBk9bRN3Si4y015K6SUc+PpXgxQip6MsytSrzLjoUxBf9oJF4CK5Ci8h5uJe6iO1xb9oTNp4HUU
+1H3jWIIoKbwenWVAynGkky7dKXLXTDz0zDHnNJcsI1mq2Q/c5lg3k8sMDaN2z88UiNHDfL/mhgO
q+sIpVUnCU35Zrc1Y4LRpT8kXT5EKzNTdKuWqzlMPRONgYnf9CqjJ4FEBqZckHUQf5RYiqqF1Uqj
SLDNmyTL/ysJmtxk/Vw3O6ldglJkprI+8Tr3qJEGAQRCYXDhxjSFehzw7SxHcegvu7mfUVntJB4I
jjJPWt383QT43SplOtB+Mnt2E5gG+gpPCN2nueJ15uJ1RFmME9PlOFnJpGadrCKQqZJDHyMNpYOf
6NgV/67TDF5+pD8if3JxxJ9e1xa5QWnkLZFm5oz8EC+kLwFTW//SHjW9ODK9r/ZXyOn8rKvEsl33
1wCtv0thrI+4FuEn5ThW7AfCyqpi2Osbn4Au5tsZafshq9mUPphGWgLExx/SQDV5nEOnv23325JF
Rifgf4U+DF0KK2X8vLw5SI76EbwBF9swxKbvTKeWTnHrikJlFvpgiNfEJ5CmMm01/ASHmKgFY/PS
GnjbLOY4JMaZ/jFpvF05X0WX4LMIpOgfjx1M38CH296/o4DoSS6Y5khVpjiXYPGs4DXRw5LKNbRg
aMiFWgjfFUPDqlXfa2AMli/yBPwAx2XPx5qXWGRBbObI+8MH4X7zZmdmmow9fB1x5OhLa53Mn7hZ
K0nNXYM9hjhUsjsKiw9/VYic8RGqPa4ReN38WcDQWmWPBf3AU7ENipkaWgfOzRBWQPS3Ij9fwd28
5bmVR8GGobm32cseKdE56/ATKcdtHAO+fvT1F0ODfOI2WYOurBvbP+jmTPKWtnAFv4XA2Yrlzno9
Ice2IK64uhDRK6jVQmOlo+CDPW5IS8Az20FEf2+V/XUZyA9L6Qsnz1EpOEQLtJ6JOjOdz2jwCD/v
iNWMEzbleZcAW2DwYLXc/CsVmeXEKEgRoaHal6lZItmewV4TTfGgpOA14zVjTiamMitdDzli52aU
aYEBgvQpTg/mVdLvfbtf2cM5YzyH4PA14Tneq6Cj/x4Yc+RaalLQ8O523672IjSsdWRRdkabUxDq
cXBHtcMSMx74XpXYE/6trgD6P7iVU3HYF35SNbAF6yPKdb8kQVEdFjMHvAGKyjnqGte2GDIqfktC
SD+s7A7WznWsJUnrEJZLOz6S9cNKp9AZWcOx4Pn6IlCuHrlLNR8QhdJLrb0vJSSAlWpFCkzxfTNf
zFEeJf3CPoo63AOSRk1Z9SDd+XsjLIU3LC/6KU4QGjQrljNC16b6ZSWC8YT2vDC9EiAcwsKhdZg5
48eT9sSL/7rnINpj9fuZWOp/AVr2Sd6zOrJmZMW4snIQ568+WWmeSpDlTXhfufBwT3Im/GNLSxxh
T3Ra3j/DuTWeVXvDEtfgLO6zklIgKMKeOjMsb6AJX+Id7OyCaWV3xhh+SwsfcTifxg24liYLAr2E
WTZaHldClfKIekQlmn5IihTTIE5nUra2WN/gP7RvFzL/kJwjytvBjeEmMS1UX4AXHT4z/TmUNoO4
z2D5FhCr3EJaJCGGu3x6D21+GftRDWW6pfmS9jlT74ImNxkMxGqw1sIiC5gNtfINruqv65Ind3jG
3Z3bGYgxb6roJqmT8Uz4IrpUkSuz/nVw3JPRUDkwNbGOKp3dZcMPd/HhXh8LysOtsEbLxFhRFWm7
5m9LRcGKaZcFdjKav+ZZNK8DXZNja7DbH06j+U2clTxcFn7DgsIGdomGVqzuFIGgnQHbkTmWoDdI
A3vjqtpmR4re/kcVJ2O9Hf7RBsYDZNL7COgyut2drHPf1Mgzi260B03/HlloFPsKjCQS+H2DVETp
gePreB8BJ82UKMMjxuKRgNaEceV90y9Tya/0NFUOCkDCUxS8d1LF8omx0u+99b2h59waoyg/CceP
yPi4xv8VMPtusq3As/7q9yNrX2ZNgogUfZU1GjQGV9Hma4qwuRktFUSzyEudHt23wZiYFIcokjej
k5cUDFxoIVWeRCUb1xwyp4FE3KV5HFqb50XJs8ApLyDmmC+gPwxJwjcewkmi/G71aEqjGXPjD+Mi
Z+xgKhqA0hOxUa2yN9ZTGreuxcTYgbY5X3d2UO89ZXGKl9ounHczfwUYib3CLTW9sIRA/AJh6kPl
383lvCpodJpPYwMSlI0uVrtf5DKMOZldIWdh746Ypl7qd+SAl7q8KE86D+YH4te44lWy6VOhNFUb
HVcO6B8Xy2Tk7tg9Vs+ufgcI3tHTvy4LXHrmbikBUae27ebRKiDkFRxV7ruaCt9TXm+S4MvmDlfN
BhEI8BmV5KkqXqzeHYFM8rWQlkNC84hemdcXiFLpqDLl/U9eGz7FmG1KzyE4/5aduGkKwuAzinIV
q5ld6BBROlNGSbDvq+xpgTxZEXH6rbWPXi96qd4yB6gw1pWJMXrv3ijhmV15LyS4loi9n8pAmqJX
fMyzlwskUG0ZjPztlyfaGdpkrDv0lAs8GfG3lFQzaofbLGs1Fhkjj2hI8tgMBpboFxB5SAJ9PM8L
cO8c9n1e9JL5RtJE5iktmRJK31qI0rhVEY1mZAc7vlC9+PCqt0oGP3rbGGdD/GUwkX7CkEmgu7Ze
W62euoTUsdwIXG0syW/uDzHqADYmnwnWcGij6MKUKmkiuqse0WlLTtkSsRHh6GR3ZeE74pkGPlIg
T1H+q95jnIs2UQqJHXgwF+a58mN7U1akMpfliWfB5HSI6/3c3KqeBeW3Mpi8DF//3nMBMwQJyWYD
23wy31ixqo38E99UNRPghiTIC2U4obiShzbrXNjnLR2i/Y0x68ex2Kbpn8UdgOtZ5XoKH8/h/lsh
BB6oNqavO7BwoTytyskxnXSAPD3gphrDMgCF/rtrlibMEQph3O7dkSDi3D5jzFMWOVd7ydLfeI+e
AdfoAQarXF5afLgrRtDSyZHJnp7rkdHIEJE3Yl0wjmfy5UX5skwSpF7jNWztkMUq+Fo/a4qcSre0
31QID07BSbjCYhG4Lbk24WinBGTeT8dH6irl/mEnPVWBeGqO4hzsjt0vc76gh0y3GNyo8mlJHpKg
IbdnqwRLwFJ9rY/W4GwpIdkJ+NZcu98DDqM6dZKzvXQyK94SuU8c2pUhSdvGdWLoQaoDiAaEAuq6
isd/3EWrNT4QFBt9A3cMCtTYkayM9GD0AM32QFIri80ZlMvPQSm+YXnSDOhkJ7wXshzsRZMW8Csf
4UIAnIIRbnUyv+p6hWtassRLJmbDnZPQpUfOVOyFontBHU8oPU22TL3kTBo1HUCL2mRS9prbESoi
d15LVDa1OASCvGo7NMejnVG2mmSjMr8Zde22dIgbqN55KyW96E2yl0ZVKBUHA5v2rrrUVwPGwnxe
NPyt5i0M7/9N7pZoX/kLxdq6ZzSQcBU4kyvlbqbk0R55RMGaDzkxZNaNwtO7OYzHgkcjvWAgKVWk
mojRPDr3bEGmK2JEkYDyPz9fRK7mGqPYwre77PZOpj8mYllJETcZlC4jq1E4UcAPvGJuvNzdzqBh
m4umiSRPTcB4+E9p2qJxVBcjMqqw/PXBY48ooKGTmpLSrFgU7Ho4Cc2ocSla32Sx7bP6U6xK5yl/
a1Yn7MZU0+Iq7UVyEFELg8nbgg/ssiH6giMJW5gXtVL9973qbLwN184VWyvnFMUbdIDgJyzjDDjm
yE94dudsQ4iZQ49f9vsY9OcGyrpTB3zxcqREEoH+ZmnxJpLBrBdodFmN2Hv5dxgUb265n5Zqik1r
8Uuhr2uUBevWENfcMsoL0cQvqCp53bqOhqAQTWFM/RI48hYjwmXc4pMLKNSI/eyxEG8ZdRQ4NLpd
J0G28iIZP9SVPR2o9KEtrnrVDtsBV68o7v21hz0TuEbA0z5G/P6OWtCyB6hLt6ePN0zqRKK43ssN
Jeef98T052hialTEtiHzY9nFfGcJATXYi6ETeB7tmpAPgTZioA0hgHzueSereORRikz60t6UwMER
jQUAsnPj05vcGpYW6mzbts3XdVubxPWmrVoTkhys/fK/HYGu1WrgrrEd+Ei4GyLSbuBL7bHADCNc
rqiR/v63tJ1l49PLocZ7HFiVIyaVEV9+eGifVb29UEUEvj0jYiBe76AWu4yTd/lpasr8L3e8ISL5
DS70jRlhq7+wavoI7fQFXAsmXn7D44pmyRqa1K0hSzO0Wr73lQdA2DoqXuMjjrkYRdPYMLQkV4w8
s4jzYocSVjQei35m2M6w3ul/QQfuOJg1NOgrFIclM0H/+aeyDt0/UWCvJc8LS+wT8Iv/YQ2pqkzS
6EUIi/xw01gi/CCdKWke+OVbq+dixaP4hJTXcLtG23qCX4HPemt1eW7W4EtNNAAWwBRkC4KthFhL
lKVJ5E45lB1rSxT7ba4qFc24r6J7JBzOKujP8PIo4I4ABEaM1sDdJGcFI+fJVnoVHg99Tc4O2mLq
gxeMh9XzC2nEuJ/A8yW+dD2EI5D4vtzZwN5BTUxIUJL7c3KvlXJKvYuBYeMQ4sCAtZPV0G1ELtrL
+ly+q1uEsrJDFkBKi8ppzLe75B2U1WElMCD8GYiDLOxl68LnUOYJTpSREtwgzkXcr+TDSfs7MtD4
8iYuLVBlpydIFExhLEfwLFTFxY9Rx6mLE/DGuDZbImceQnMtTH/yR/MR5QCAD+Ameuaerb3O7awD
bY3n/YNfki2T9qkN/yOYZnT/AkrrddmIVLEGG++pSQqY1diBe8D3qQV/evJB7WQqKYQ6zfBLZWbi
n9e2qgDVuPxhEqEYyBOpcl2BXKX7pr3HkOosG68P3xlUKJwgCLCuQviTzQ2q1e4x5mAlv8+0IGcN
n9OF4rutWQTIgx0DV2D/ci3SeBMVepbeOiSiRyS3XTK1hDpiY9g43d+yP76YeQA7vld79Pjob48G
RWft28TqfOREtdgMfmwo6EQwD/adoc6J7HJuPYD4hoMzZXdseCrzk5pYIQXa0IgoTEAvifc3Bev/
TgdPrBg5ADmC5GysK0KLYDXNmYSbVL39hXIPjSnhheeIibeZjw50/YfPWRxHCL+4SYh0k45KBlIl
IeStXz+xv4PB6FKZ2o7ckFqZvulCR5Ggmi5xAGaZuh07gz+P0mFW94V1kdJmSye1sZKca713ILOh
8kxvm7s0IEvzxxGyFK6BuxF2coamqGWBvHZ+Gq37N2QvpV/bm9GTzsZqimxChVPTks2sx+dbqH9N
XGgLW9B5AdvEsNdWJ/s9kKPDBjP3gf08CNqDVNFu6oyCrTr71IL7IoCI5sSxl8Hhwd56OHFzQLWC
RF+mkInZAQWwk4zdcW+yM9Y8ym16+AOG3PfTkBOV/x0H484nxIuzBApLx8A2IL3SRRFelxkSDEKL
UHQvVDU1j2u5RwOuTzYhop9dzqgKilixTgQaoAfzdjAl29dGsU4AHuUp/ps+mUuPbI0L1RxeZyWw
jxtr/BfFPWD0igXlLD4vG+eoxAsnvM2kTG2UuqaEWozb5Kl88sUPmvPJ08ANASvHcq/qkDfIAKLF
MrdWIFH9fnJ1EmKZwGpk60vIaJWURtCnb+ejJ6uoJQZ+PPWlrzENgYBCUYxKT2ikN7rPf2aJy/lq
q5442D8CWxojAu/sthVsHlkUpX+cKtljXp9y6Oz008BmXX1qKvITbPOoG3DBwraA0x9EgscHq8Kf
LkFdkpzA76pBXa10x+iqOQpsEWS9oywTx20ef7PcmfgJVl9PWRrs3UxbR7dSA8G87PLgDoN2F/aA
IyCOztWYAJqBD1InRiLlYS+dNZu9slEEVh1Qt5rjJa6yYcezyLMrv9hln7F5T3eeFDo22+KsArF1
9LU2qOp33OYOqwQp9bqrGErEL2+xLXuaB+pgR+jGo7yBuoYOJk38atDThsAt00wHf8T1hVnE5aBf
QLK1YpRcuZg9mD9ZegBQDDgXkF8IhQr2hRHPA1nZMkVRDgn+UY4zyjMiNi3tqBOxzqT1Fg7efkqs
G65shjgZuTRFwdS9Jg6wSx/WxfFPz4Koe8dLH+SA6YljQvtTys18Hxy4yYldBg2odUoE5SQh92X5
YHqClOEslb/uNGssnOhS0+JE+UIk5ab/5zK5IWJ7vH5qX7dMCaChzoFXe/wWWT2qf+Qj1VwgcNOw
W7o42BY/QoL6mWE3A80mM6sjyKQVtiKEKeslXVxZg86eujip86zxW+ni4cOYoMr5c/QhPpMYqno/
9PsL0C0r21HvYtVCmPjVCVozrFjrSzX40t6ZYsxpkDtWl/z0mHmZTZIGieSJu79G4OQms3Lemsu8
2Z8Ixc2ZK7u6LJ+C01HJA6wvHwb5j14Ult0pf+VkVyB7c0k3ll1GIV7B7+wC9M6u7KquvAUtVE80
rf+x8c0VfDjW8ux16+Wna2ZBuw6MeSgX6AiFQtOrEiihnno/QQMlak3ssEBIQiyBa4wJQGyrZhPP
mQpWiPWE23/wVsubv1GHjlCA+svw1t1HZZ4n8Q321aUPChviemlDuy1J2z67yvL4SbAZENO41zzL
9WkdA26Q8L/GwBJD0981KXnxuirPlRE/u/CAMQV/+cIDxwQvJvxHiC5pxChGg6OFK/eGsTNMsTsX
HY94KOcF8OMhU5SJcbhaNoteP8ID7KvmJapgG+dtohuzIQwzr+FntB42RYfRmYy61TDYi019mt2I
HCrlq0XC8HuPoSm1BCB9v0M6XicSVNHMBsH9Am8R7z7ojSJsbCntQPOvnbbLjRrP/aorPqJCU7Cp
axDlP9vNf7LoCR37AiN2z4c4BfI89GAK76RmRdvoronOOE2CtT6SjXI3QgOMwHPofm/q1ve0SQVj
ZvCqzSAtp9v38Khzz6HppSHr10zbD+zWpYH1b8dNuX6/4GN4MOLy7uy8C3QV47xp+hmv2yMJS1xr
K71p8dto+1MS1DzZ497GZdL9FK2CwyjNzPwXjgb/GVRklF9YdzbdNCxm67YPJt4GX11aEbqBbfIY
uieQ+K38539yV7Fyg7AuErxfF2p565N9rCKXXVRUy3fZLfjnWxqQ/7kTVewqgheYnD8HePg/xpaQ
uNEgEnaF3FEZhxbtn4MZUqwwaF2zdh1v0CFpwQuP5qPW3Avf24Z6CZWNR/trA5fRru3u6WhGNang
AnVCYKpFyIn4gCxPVmdG1iUaqCCPXsXP+jM736D9yTti5oV7BMgNzZqjrzFFPl3bnPMFdh51m87+
YTEcC5geQkqG/0GXBEK+3UVjFyd/V89yVFZ8G7EoQiP5aZBExBvlMTuVZDeiGfsPsoZv/iS2s8HU
pJXpePJdxBSUbVgKL0Qlx82dqh6lApCa4qGDWfvwqXquIiL6/l/mTiP4Kg5G26QluC+O7AZpKT/U
/f+drO3dBKhRrEYxJDWYxOl1gNjq4X1uyqf/HT1HFiDJKkvR25tF0YnJq7yuaBwFi5Qr/p1b8NjO
ShHdDV2KZJ9Lk/InzQ+E5z7Y6x5IRTP67PlvLHOZayxkF4Fm9FibyZTrVKcqSK0FLQJwEqk/nw27
I7wX9mXBmMBJGcIDB4arKBtu2fPUtTWTTrWFyynI1vauH4rhSPAN6htJ4JoTwcwxGr48K2/4ogDo
O2V9uSSiponjueRFdrlXIENnhyKajjEn1stZLso1fh33iVsIMGHoUO7gEWpdpDU/pC39L3Cr4EEf
8oXQA7Z8n4nXPJ3QLspIz4V+dcwe/qiIkYVccA74mqpTwT74VWmu6syjX4vJs8olCTsVpVlZFUAq
E+ou4fS+pdXE9l9xZaYAJl12/JP6hbKQTtrsXC9nH5JMlgtTSB1P+ZTJ2PXBnoUjXj5AYXrHvTuV
GaQNYjmDajKAbFRoUoJeKW/qtwhoXXkpIAWs7c9TMn5Y0GP27LA9zyazj4gRh4Fp0MSnm3kyMwWk
v0o3yoiexmPTBxuGRnSM8r80PkXay7n9nxmnEv03A0XK7yeT7HVLH2x00jcuTYFzLOc+LaEp9/hv
yab4rDhHYq2sMgnwywCt2RMVV8UkP6mfoEjl8BQkINoySRN0+pSkr+r7sF4shycHKzptAkj9doqx
zWz0wofBYuhEd9ntCqUus+i93Hhn2yaRJq/hx3erwz0ANSMgydmxLoRWVwlIyPgOEuWcMKFO/3kh
XEcWUuRlTXAUUKtdpLJ2jzNTPIDKM++BuLin6NyMoLQdL5daDMtEaQYrEx1X66qCUtKYNcLJNoP5
OmZto5PqpE0fqkLLWqFdmeGRCC7+1WnA9w6hh/Na5Z2Kx32kPq3NVCAfXqOr6Z0sUH+9lw56oamz
fDRYI9iMJG9mGZsRHWNnT9AAX+FnGAUkxY6OnsMqCvRftoQaZFyUyswLpApyjKgqE+hq/FQuJ/UT
KyFCjBiYQkkeCOCFanC8D+FrzkonxrlU2sr0UfbIs5nshNERjxSvn6KsBR7twj80n93PjHuvkyIq
IUhbHZrFXpUqxIN5UnAz8TKFxUrmeGtGOVd9lJFDkmf6dvh2rVw6xlKm7Nq6aoTjjiGLcEYXc5ut
Pg0i0hbPzlPdK/DSR83afzZPHpu+Uf9bQU/4LuGyH2dZyEE4//bKTJLSG4t8BjC562JsZd+B2RCl
BApm2Cp6EAYnejf76zghqhX/cx/yt+x/NNx1h9V8yoQ6qNrjot9qeEixk+JDnneOEbtgXfb5YUk6
gNkMzIj7rdtaQI8W8hGCXvKKAH74eXhfjDDHCoDwwbMi1xOxmi253FrxqGEexCgZx/NlDQZmXahs
441eE/3REXO4Qp5ykrf5Ziwyd/E4lQJRaaYVq5gqv/LfEiC2hYduFQPECUpIIMdApLawhVQqXAyU
VCnF4Pma34/dx4Ynycr70TKoNuCdDpv3BsZf2Wplh5RPoDZd05NSyleCAKcJgqDbC7kAd1wKw1nV
EVMns2xpICAue7L/oHZ9rzZHIgyNavwX3SUSsShVItPtmFvl4mb6OUIzd9j4DBp9dSntnoHvcclz
4KZUn7fmb+4iQj4rNQso0hBCsfs2gzRXtzcmANQDo+WnBFFxx+M9M3pGejhhcUailZlrjs/ZV1OH
QWj+0A0lSDOS0RGuKws6Jyu3zicystW7v6Ij84akw+mPFCz90lo+86IdMVU67L+wKqsHtEfAqH2b
j/1k/8xoGXApZVNxgs/+aXiMEiMriPe3/s+pgMV2iDalcMhN81nmkQobbJqMJF9EUxQVTB/0e+Kp
23i9asuMlqKdGTAZQYtS8FZ9i7rBNgdLtMUzHH7Nuj0bPf5W+z8o6V/tj9HV+CYFXJUavrnHb46B
KvpY59QH/b221rawS8fxS6YRPZ5J2qGf5mYsyzuB1d1HNexFpT0lMPysBzgkmTTjuywDHQlD3pM9
pyGenpDUsdNXg1ypdfLrwAu7E/CUtKfLFnF/myH68luJFUTE7+fP8iflnLUZwiaioCQhGQlqSIp3
TC8Zx7IfZo9NB0Ma+owogXrUxMSKK5Q1ntFgh4CcgbIe8pLVYSnb8FQiq3W7PvIM/qeJYuKotczr
5VLznNLFaGnfMhl5/rVFCovLqtvc8bvys2ZjeQtNQrbn6Y4tMCvsWQ/4i9KsSxd8SOLPitNHpSH6
J1QqFkukbck68a07ls61VhJg+Om37wWExoW1Ny3OxJ1goGFfVz413SpOl7ILfpSenxoGJBWExGAG
wbvp3ByHFe7QBsIM1TpJKCiqe+2LFJRkmVzl9VVLvkDjBC6cwNbD6u8YdyWrOUf8KjnY+4GVXiEP
Xsk1GTnystmMkS+ODdxIZZTVXjAg+UwRx2DK3jwFWZQdFZ2yv7j5qxQBh+YHzFiaelrGXH3edixJ
XoyK9Ps9n5pfXXxwRv17Z8mAYmUBdmPe4gsiAZd5M/Pu+7fvm1wc6iTYZ7udEFtbmBEmRZwJnABe
ch2LGHj6e1tkJ+NiD8/NlAellWFiapQhZGEiVWY/8d6xsNVYcsDd+D/N/O1Bg9/ZOGSR1vgdnv/Z
iJ214uRqvrpWzK4dD2yV16nanKepEUstXNq+Kaur+FnwNftFt6GsOexznCcGOoFRc43y5kG/rjGN
6D8DaXKZRJA7Qk/ULeJmSKK9nWJmSoFM1ATewytmPXoAe7cjB4IIauNeDNkxbbeNVT6e31lw3D1+
65Er/sFlzDbfetaWr4/plUwobMOAIV5D3lrWgLRu/pff8eiU4uyjn1kamwrWmm8VeMiImaAJtlaa
bSYxUqG76mXfMceLssLkrdAPRr8kfBHg3iZNpnrQnAxhHhwBaVWDv8I7dcETnPi9aBlrFLhcjMoD
muAFidZYzWIo2yyYC1qjPbTi9C33ZOhhOSRAJeRJEixglw1bX0u9i3N/ExnTk4XAoOlXYdpOjMQ8
bKpHHWFFGM1/IVDx1KEVJt0SrrgFA1CKXy+N+/GEk12/YXoIAydCztnyq4BFCdR2vUThcTqfP/9o
r9FATSJliwZKgYP0oO7QDpS/EGO8uMihAyx/1HarU2u4x7SV5uyFZEbed+qpMR1lIpXTmyZQ6alO
s8KN1BoZu0832Ts8mkoBa1A1l4g3eaxTWcxHpvKt7stSpLPTCGF8FIN19qXQzZjK7Vv1jOf1Cq7l
eL+WePdpbKvNc/+IijmrTVznRp7fIM2PIpKPWIa0310rJrxpwiCK4I7KKLm42vbCALYqpLobrpYH
D7ZxmczZrH8nfdxXK1yzL5JzOqxZN/wKJ9WYyn2GpqF3Sh19Gkke5aZOxtjMP3wgW56xwfVwgO27
7BM9b9QxJcmAkkfeyQBGvrxv3AnUS4abkCzujHCh5gEFSgj9+7wboqxXUHHiD51upYlg3Jlhqan1
coKrlBf/5uGPdoQ7/+OqEBJXsuPTHoxyaZ9EiA67XfiEtMSDj0ztpORpQS0+/tLMp+DBCum+J0Qo
VZ9FQcaS52IgS7jmZPtliFwZ/Ccy2/qpjXb5fW4c5dX8q0XWlI6PX4RTPbRk8Usn3Fwyrq906WAu
qsbqyFcU2dXbgRJjzchE0irPRQREn/2kO2gODzOQUbghazh79acEvaVaRRNX+oSbN9aKDQJaD6Iy
yXw9d/2XJOQhl+9j9v3owjW1UJZFFmBMVT3qFXfqjUHPuWQvzNK3RBXdObIwdlYqZHm38wjAfNso
G8TAz39+uWHU+ss9OCjLnfUjjqNhO+0nGBlB465UZLjnK9CpMWzA5NNudRRj2fZhZK5ueIY73kpR
Qi7v1GbRZQuilDRHH2VMr+LuFm2Q3Bbf3nHi6amaOGwkGNahVuWtd+xm5z/ywlWlYfkqxHLOy7hp
3d/G8YlaWuNIzvxw2T8HELJZmtxYw/q6e0gs1YpZngl4+XuM6zE6EGDzPqGd+dwk5p1NlshfaL8H
cAvTGewi3wX9+iCthOCKKc1lytM++ezLhyyD5uiJb2Ba1AwNuTo5RYQt95Tn69rO0ROmQaYLuSrx
wbvWfz/qMKBI2igT3b/wxvqazguWCnx3Mp0pjSZmAqA2Ak17Yd56OxR420SEsWws4tUBeSGPsuXL
Rw9PTphNC63lQw8tkHzzRJr907IEjNOCSH6DR7Z7EldtgoTPNX0YkHFKbwP6jExiW6IKtV2Cocwh
08nnN/XozEJc6JdAtFK7poS4r9qpNwJIwoRXZpA2VRdNQp9QNYyJR2W9FEmqBLNjydPBR+IgohZm
QlKPGu0lzqfPlRuz6KyyR2CTKmD2jkkfB7sphMJ236WPJYlTKnDz65bxbCFkb4NkAOPYpQf4RHCb
XeFhaLHmtOvUf52xV16eoUsxWWlpEQKSlvgFkRHKI77vTWxJoMxDAuA4MWQYWYA7YW6Lyf01yxJP
3Lojf2j+XTUqu24F/H5vAoGuvWA9jDK958bwtatNzDRbeZZ6ahlYJZ+8JRnSgWjeMuwp8h3gxLIR
570xDBl2IIss2oCXcXutodScqsrX7eqMPcjZbY2ZJqc5nZGfDtdM8M8kMHeobsnqKh7B16vOj7nd
7gErLvuRS9pyTA6IeQMHTD0gkfCLyi/8x24L0Eh+SI1LIpc/S40Z8tzT/UHgQPmVPEBU58Oz2oYk
DMi41a7CZuInH1eb9ss6rHfDAhvHbXyadIIeeznc7X3PbyZaReod1PDDy560WCfGpSEjQsl7SgJk
x0lghJhpxkTOC09rKhR2klDxYSAkhvfgGg3tNsPcNmA5jkP/6xC3wCA7C5N2oLiu5R7TEyEuzp+1
k1kE3QsNLD1bYJCgjCbvirSPiEJa2pg6nHW3bmUzSeHt/tO/0ISEWQr1Nz9u8wSBpmCiJHEPdN1F
TRlfT6BLzH22n/bm9hsXPth4vE6HIkwlJOCQyGp+jHmgZb+bbBGYliQPYX4mrpUoQSr1dE7xiMxY
Y56TsRapw4DUuecLTb/fenQ/Oz/B38tlZgo3NH2PpUDN74z6LM1Ut76Jyyfl+2f9LiX5OARacLf2
2+ehyLh5zw6dUYgYPmMmLl4jd0IjN44p9Jnb8TISF2SufzR6gtGuvHpQ749Czm38pU00BwHdYCeX
I1Su5HOnq4RpQ2kklx50qvBjTX7XV3eafw8v3Xyj6p/ALiGLSkHfyXX/yTy+7irBphHXl36Dbyv5
AsOLbQc596IVymAGgN5pIaxrmiT6+lYFI7BkmlkcL+QiAiqYqACNnJvYRoBJljXQWkCagPBgInup
C1XbtDJPp9+9td/eCuqGJ2s5/53qRw+CMyxkBGts6sTFcRiS2H+d8RH13YJNDnsssiGxXX6LdfuO
+tmCkDNHW7Eco4NHOzkZMSZ5kfNnrKpZ174SSGjC3WXOhG+jwuOtqJ3Dlx1LxJtebRXjkINyTzM9
afvuZKaQPgjektD9duh2AzYlltodpwcDLS5BiCh4pUe03XWyOJPZb6PlnKE+0ETNaeneJQ9EqBCQ
vC0RBIZ/ydn0/G1Ljs9khoPiGZr5V6T4LQh06QSDO3YmHbbYNMLw2MNKoyjn75g0bsKv3kxsl/kJ
bZ9TvbMeYeNcf0BMqynZ+fyFYhiXirZ+7wNlLwjt376TRhENcjKY/7/OCAjlVlF0NjzRLcXrbB66
hkyHID4P9x3HdvzRJTgQeA3PWGqXT2UpB7wiwM5lRla5BcHotwkR2PQPiSpF1thSj9e1tgWuxHUN
Om6fvBMKjhfwxDK8k3ZSJ+R1V3cvLx6svBcKRGnl9jMMLNmnAC0ySiDYL5rQM5cfvy+9ey9oc1pn
lDBRZiP7T422OW3U9YqUkGZvOhu7JXU2A7Z9iYT0cUgqgwnwxjNLTsZK0DwS6mA2Cy+ZFqVUmtKk
dSz68n0b8VQUIPqJifkj1I5FKiImHC0t0mU8m3KBafADghuyVlXSfKzRAEDqwFBlgu0jsKT4uV3v
NwAcN2IxUPHcNcTGWwXtWoBMMVNb9NvoMEzmWKRK935uJAsk/GtRZ2ih2vowtjWksn9ypZmLjhDA
vCQLElMYIb8lXseOJBp5MoRBN006eVaxe9p8lg4FeaQdkBUHvQJZxr8D8vHcYbuG8j27iQrv2DxX
b6f46ylyIWS8SvTNFOrowbg7bUaonsqECrbckQ/FSSsmacTKlWo/B6ekisdYt9oGRlnMIcTMTccj
OEDfKUJ9ZTxMggoyIiI7vkyTNTxrpRBlv/FaoVXVvrVXuHgLiQh6bhrYz++QiTIytv4NEHwWYZ2e
ah4MZ6M5VCar/k5UkPDM60lLcc3hsMMhS4CVG+p8Ld+4us8OowFQDrx7RyD5Egx15TsTdo+7ZBGq
7NP4Cyk84NcSVV5SUVwHf3Ip4qg7JmQh0PqjS2YT+3AWNgR7RD2uzqwsfyglEiKHdOED9dnR9Qia
TPMuS9ZOjbzdIPV7xfDg7roPTK0MPrdRGJGhKQON4PTevGA9gorUsEqTIU0xk4pDMDA/2w+3ooUx
5u4TRL4iX0sr+dt7W+e4bhkz4XDKvKUVKdqHfgDeZgfeKcDgWSyQBJLG+qGibkAPk2ZYYNEinmuM
XQHaH/pOKW7ASqF/rZ4AwvOPqVEECeWS2AFSzyZO6PBn+Y174pKUEy433yKqYoXnHq3TsEsPwtm3
1ksJRkE888EQA7ZgaY5e2bw6vrGXxzJK4Cqae/VxFIIcN9/fI75H5PlyAkclLG+59pBj5bLiUDgW
jbFFGJpWIfPIX+3ZZVHNe97O3i12UwGZtPzD7cxR73ARvZbYagGq9AQAP7fVn7iC4sE88pSym7EW
IZzYgcm9zccnMZDED+r3a/SRccJZ2QesCcaEStpQQW90lch22I7yzZpP+aCNotbtse9sIIRy2yWE
hHdhFIN2HpCqy487Gdw+MyPyFIVUQfR9fyAWDStU+wQMHi0hTrqNFBKE8VU7M9d+gwNsqh6BBe7W
z9vzXPRswDbfK509s0IJ4eV2UAtEQ2L5ycSAtIJyYfsDbIp5t+uP1SB3l6iZzflVqtHlEaC4FZ9Z
iWk8uMY6wAFhalNBHgSu/3PAMY4gxrZAjC3Iy+W3F12ikHcuOWbQm/944CNQA/0mnUvgSAPGzbxg
y/OQz6l2Y1ypby0+IRavJKlsY168JE0klpvErmWbDfLmDA8KtR4ntp3NtGgRrdaSsg62DRLzfr3L
YIxzlx1SKHbsXF/zpeKOmdUSEAapr0pPtyuiyWjh1R63mzuWDCmpXg1ALwT6Q/HGQlDLGKtiOFHA
aB9244WJcUotCBLQZe4RFfYLYxzl47GVpe9fx1qk67rfmgqCB2ZZY6V9GiJSRBUZkBB3uimsDskV
8mtjrWHXjJLrava0l70ggmUYWisebuCoJkX3NMPvpHpAGYheqsgJlaqvpE9yQ/SfgEOgY2gp2sc4
SMFpfsTJj7tAXlP144syaeBtZejg2Wf3XtGD8YcnPnoU0U1TuRBsLSB2+RBn5mr6FJ58r/ru+INy
UZkL6Gy4VB4PdFZXJnK8iTncSAnew9M1foemqHbCAsF7F1wnvYPCPqj2+cg23F9RUJpejwnvnBBQ
W6mLpqaX/0PQscuxGlR2RWdBUM9x9316cB/OM2WDAUW42yd4gRd9qqI1s4vfccKZuEn54qRhZexR
grlovasjtEtqmjAwkWuaOHlpoWWyU8N1xo8sOKTycaS7hJEVIxSLYg4AwvGRayZnDQAc0/62IFUP
7Dwr2fMeatc0lsK0woJ4qcX6wmkqFCkFxOllKB4lR9VoTgFdt2ANRl4FXBQ8eYGWf6knf2dQaNtL
a57+fuzrDtTuiUuL3G/JJdzFY1tpoIY4dHn/GFUoDTJZ6tM5dyz3Yy1WqODUClYlaaP9xRQ+HGy1
JwlTfAFsao55q9IZMeRimAotqIgrXccb53znIUTWc9bWbI6EbiGGVwf+7aRjQ4qnJDpJAnjQZjy2
VigUzMve9V2j6qbkotMDtCBBErozI65IbRVbgVgEEu346JdeId0QqJUKuN40HkXtDTadCYLHwvwL
tkLMcAhUz+X7se3piUOeXvS1Nv3VHDlTYGnge7xcN4RUD0M3/wkXVTQk9+K9c+1cSZ17sIyhQtRs
9Lnso5N3yzj5oyE5QS4pNTqc3iPSMxwv9FUrsJLC2JnQwkVpdvJFDKWWN76qqbioUr5bDGc+YHJE
bhYOjOp2jsnTRUXbcO09zgWRgBMTdzJGENOAxvwaq8oY+C2AnKu8XE/MJ2hm0Ppi5PKVCEJ4hgp1
MNfOggbOhOmsXg8YDDAx3lM8GqKTCKgc392dTW6LlUJNM04uaxKOKjnq3rXOnVdhPeliwN+67MYp
oQhbSoKj6I0r2Vh4JCpQ0dEM2nYwuDeE4Ag84P5T+9t8TgqdZrfyShblbkB/IVZI+RPZ+bK+7jGu
/J2n+UqHUChcz1Ab7cKP8iSBxvXYo2uR++P/BIQaccon2HXTlsqIrCMU0kGKL+W4sYvaAISPTL6/
uoAZmPHbo4Re5kEhbK+3cYKN3tdkdpDXTxnYEtmb22PDU46WoiU8OdRSpzz96AdMBrxeCBj/MAib
gq7czmo0//y0uZiXky9LGHOKxFMIQ/WigGwKo7WLI5IXvmStkGeZUfT8TZ9bv9Kbbp06qdPkXJax
3o5KrrMM7/KP9nLC1ES/4cJ1ZycPPjOi48oRGIp/fQmEXal6r27Bg6r//npBgHeAfaY7Y5gQetYw
G4elmf+k4qe1GW2UXNfye/6SyxqzAUy4HSWacp1ODb0o2v8YUBxi1CJMBMwah890A+7XYki2Oc/p
zVL5fqjPunrd7c6cN0U9eJAKxNK6gn1BPvwJIeGMtEO8dx+hOOiYyUrQYaYic7FtXsyIv/QR8WAc
C662/e7ws3QJ7nXmPkol8HV6pIkDslPBM0XkhFprJQvSFUZAwuQs0gG07DCiQZts7EzqiGyOC2+j
RRPs70ftv+riS1lEb9p4G7cx82inIw0+RfYhJfpRiL3mx+zEJMPE8nVU2In8UaxdzhlaM/sZeP6w
IawcLoWwFW+/7eTQxqzfU3ZhOj/4KsOd5trcsF0TN3zMVxVdoARVNWUPE/mpIxP/BKiSjGYH97f2
Ha3Sbkst6wvfuPe7hVkjMrseuYpW7V/FjVQY8SX0RK+vJbrghfSWBs8/yUrU+uQsGrlWQlIgg1vE
xyfDn2zd/8nkkJ55fXgwZuYKBZtkJkpiJAh/483uwK6ScX/GGXkEt+25UKk5Qya7ZsBMm5WwmBPT
HU2UdT8lEvlvjFcmY0d1X1zjLXKk4AD6xW0CyMI9xV4l/QpH2ER985Pu0YGCC24hBdlyE3FE3K8v
2sKgcO58lz2hrrGWlNA8rJ0XYaJkzpXVCOyDu0agkBi83eH+PrqWQ8VRNmjDOH7xkD8Zpha6J3wZ
PzO0udLrtExIEh0MLkbRjZ7T5d8JbK5nLvpbmEYcplThbRgAya7f+V8WJhcBymtGepN0UGbL/1HZ
XuL4Rna+RGR4gNL9RdDphdL70OVaGCmPTSllcQFO8b2/Z/f2SD80U1Yf0uq3HA+P3aAOFpnbvuih
Y1SB2LoKeJiUP/UBdRZJujep0OfjO1gRjklk6YOs0ECupUhPJDtvUyWvbxyiSuE0lnbQZB0sCFOh
zIPHKLCeXI2Thlys4QB85iBR3WtvazGbDNS5Mm9COeyLeP2xeODYb6k3PNYRaLBcRSidhMb8Jakg
9ppPijTPa/XG3mt/QmkvPo5dqkeYeF/k2XPuSHxcK2Iim49tJfWrj3rctCP5PYH8iNILAoGvtIt5
y03ISVnMrHt7XGKQIK0eQLhA/FX75oos4IHMYdI3+ebEWV6sR3Dl5e4Butz5un93q/jL21OulliD
vX+JxzXlAhl5kiTC6ncn0BCAjROR5sOrVsEYQN2vkERXMBwzdMKJD3c1zMRwzrgmyyVVMLvXC9Uo
XyU307jTcneayBYNRMjp8/RJyOZVaLRTSak0OwJ/lhCS49w4ouQWC5EjN5c9kbYu5YZ7hn0xDdDj
Iobkg5FownArAyqBBFlWuvT24mtMexTddQV7bwraW7j4TanVGFeEEeB8HyUx5nlltWCtd7CGYN1c
SiiMKPqIzRMqnpGPMTcnHjSJyIgdjn9l3RyOJlvkV5xEqf5d/wwKt7QKQozxCvbgAVfqEVfp8KgN
mPjsvn3kVIZE7yN5vdN0LH/LMMEZ/faWdrxdhRtJTrBiF4nmAKBuu7FY7EaodYODpOInMmSKmcCC
Unt3i0xwmcMCCtNYT4XWlgFOmxJ1MDlgEbTr3tsWzUYGMTbnaFVeoaXHp5xOOk6KmaSh9TwMmW9a
thhkpaRRySRUmjqeuItXRf0+9KdZeAmBT4n6M31pd5stRAmk31zkmUSFSodlIVE9/moKBRw8dG4D
8MZser2LLfytVFMvIE9V7sK9KdCNIJryOI5dDfi2g3NkRbU3N69Zx9bPjOnJcVC2ELF20ujdR0uH
T6ufDbwkJF+YqFKsBiEMfiKWmeDi9eIuwCY736UID2LquxbVeSXhJeny7YQiWPnHZc+GpyRYc7ZQ
WZT9jj3C0usEYibBKqJVFV09PC4NP8oSIz33aCIt5aAIr4vtAX0ZxwkfqePl8uE6PQ7cgfxCLs4C
p4vqnIJWZfrOFGFhWjEZZteYhHZdzpk1Rw489CIZq3z/o37dYUC3hG1Ma6h/5dj89ymyUIWB6pQb
5/6Bus402hCsrO0rSNpTHi1pdeLdrfN2JQP1EDOrxTwq3RjIwgLEA/pR66BKswaJ1+o7bR6eyTbh
6AMMfSMN2QDUy8pgaAmfTVdfrEB5hoWrIuSIvNd3HE/rMPWk42Jb0a+vYIgQuVGH4Aix7LgqH1gr
BHPKwOE5ULVAFISqgtKcSIMBxaZgDOMLQpgs2X8mK9LtWJpOrW5Okb1h557KExUjbO1mMETm5ZMm
ctVS45jGdi9jEi3DUnoxLv3i6AJR0DMXgMxzu8KpuS5AtRwYzUezS3vTT/UUZNAfUjFO57m+Ij8u
KGPlWqbH5gdk6iu9SaXy2FeqmJGsvMmIJsLbHRnysqoV5eM7z+eqktgAHQAhIOr5teYNSKxsNjhb
YNJ+RB6Vcx9QhfrHLMFbvJhR9awFs5Q8i+bE6FV5ygagUnQzIN5WTmOyYl8hTYl97wu2oEFwMyIo
DO/Y20RU5B+TxnsVhRBzq+AJBbUWScbVXwil7at8HW2iEgPZokAL/h7x5tCOtS7gmcHtnTocLIl3
ybTBsAomxC/TYA/lHVz6itCaTb7df9T7t6zSwvOGq/yXVA/3i5PmxuL5hjvHR/dXiMDAykaOMUBK
3tKmUvwzuLQNThpuBBwDbKGB3En3hsgu0QaVOHy0Cza2Q0x760RTlOFiAc+7izmhUJjpw7K7WOSN
QIsW7v82UpGpJmWHBFeVxjKj/dQXv7VjoH3dFLdLgFPu1j84RwMxHxtJ1FTszEOtoRIkK/CGVGRp
rLPBQGJTYTQIkWWS99q8xoIZo2ygANl1EPAv2TyacqZBWBFFtbnAL7Q/JWpYOYAD91c3B9gZoNfH
bohb/1/1vY/maXQ6doZpscCsSLkxYUMmQQDvmk7TO6FObTxMxghZxL9rqtYet2gYg2SgakNlIquf
rhXFrMfzf0rH1vWW/izII65NQnRkq4yrpwrW5ZHVqOzhYeZbFwW7WoPckGjopFcefxe2OAodUetQ
3cl2gPdKfwToI/QdUkqRnd7fHlvMYtiPU53KCKUZsk4OrUbh5e5cDvh9VYe2X5zawHmv1OuhKrfO
h5Cq7eI/9X0iTFqOdz7VAFUVkDL/GElehyBe8tlnBEKj1PZ+c5CWWuPdNqU3maZ4gkk8JYvjrX9m
N2JeQL0NW1Q2leG2xsp+3a/6YYuTzT+rr2Pp36m8mChxa04KcerCB/w7Uy5GbTIdn9xhJUmwxZcs
lXmCzbKXCInUq2U374znUiZLmOH4I3yY+jAfvWNc2a+j7YN1uhR74M9qIReg7jskaF3xtgyhKuBX
3XO1GhuaBzBVP7I/eqWZrKWc+0cjmUPRN/LdeQPu6quP2iEoDeILAzJSIdevQ+nOxBaZ6JLzepmF
rD2FkgvUuPx3XppXu+595/g8pu98Ou2iA4aEZ4p2t/bN3WTDtGfY2g8oXyfdZnIhEUSz2mDbGffj
kk/SFvyQYAwRP2R6lhtzb/mPszrSYbQksNZ44umPHIur1oLZyXzJKzT2m6v7+YsQIP1G4TDWMzXt
yWWjANi1fg18YnFBojCe6awc6b5SARf0xH7PmcZRepxXsIaE7Mo49UZmVxqaRtRMHDDwPslHn10e
RC8FZJ8gPCR/Apm0TAtqffpFcFGr59mf39AyIz0kN26kOmmB1irw+CKpuuc8InVZfEZCv77UBKBo
kR+C3ma2ULDBlM2KhUqwDiWnpHH9DZD8YAAboWcHCDkp7mG9JpcYYF9d+GguK/fGYG0w7fy8UFBG
7DrwQ/pxdMWrDMJw0bbKsG2B+6gAx/K1t/9rtqjed7zTU35tMu943Sr5fti1jLTymvG770GFdGFV
RUkVSzpFXaY+e/qE995XcDailuCh1MTTwF4HeNeiAzpgT1hzzqmfimcXQ4J1KnkRr7UvPvzWGsTJ
YA7YDWO7CvkShzCp8nyUnyd9/hyLoBIC/8tphDvGQZg1TALbg/nFjybzVOcrpjc1SJ+zxpVAmSzh
ND5B1uty87h3PE6eHTo/uhAjYPOIBAPELfOeiy/zJzJhper2vuxq6jXSClzWvia30nZEf3htk3dB
u4c6G56zmANu7vXxCjxAurD4xWtGIJrhHM3dFiOswDWstRbYpFDjblk796eirxicgHkbQ4KYFkQi
khrxg3q5kbp2o4iulwegQTNoZrVo4QXILBtCeTrLYZI/hlNJhX6pkeGtfOgWV1LVZhnpUdjZYZP1
S9zC933H/SnI1vyZoFeI2uhyNh1HjcgXv5go2rqFj4ErUBPSwyVTUyI/yqpWJunqB8EHnGiV2lff
pA/9tSqKWgSUb9Y8iRVml/hvSJOgSMXWab195NIgF/GWXL2azOgWxTmtnIWWUwtH4eU1nS6XYKwX
GyONBdeBT9QyCPuSeZ08fVONnAW46za7z72sBaUgC3kwdeOkYdDUNKs6IsPJcyir8B/VLVOB69/I
4h6gzGMYqiuTRFp7kggFFciG1j5W4JPTGUNMllIa9BcQ0gJ1QxfJ5tD/DokUrJY0YtqipmmtmOuH
jmFjD80SFK2Iat0XsQ6tCUNzaSwSQXrmO/ITSq7iUVoRee+4SBuJ6gkYWrsJaAvfPO+1GCJGmVdb
c1fVb3yli2D0gU3QdLIR5Hp0L/7/b3id3U9Dntl6PloY8zPXHDMLMGQZ7hRbinXC/LD1WZgCkhpk
knzmZk1YoWewZl3OqzRoSYQcbaD7Dw7Ko6FPZL6paJ2hqnu45ddSPBVWkFeVRKweRndMe4lOR0Jh
+LgUAoit6rJuYC6X7t2Fs0a5lw6CNUBgR/9C/QB1UaI4yLrLVdActgTGFul9t6kCrdfpNzspyGB1
EW6NGgF989zR7w6jZQLeLO1ojF4UomllaR7OxQWHTtfSf7ZcW2FUoUa3wT6KU+xizi1O7fHxAivQ
3d2V+w81KYBvIhdPaJph735+3SKTFBpyyS37Kt4XaFzO9TvK51yBsqpCU21u52jxnXJLm1JBGmOg
7E/7tLiR2mzzNVFpX5MDkMo4tUtkmlYonZOnMyEZM93S1609vdCL7c2ZBLAwzFJnU8tvOREPAblR
MB7wkRGhoXOF2y5uq0o+QempWFJCa0fUfKHGNRID8fUDN3eah4zLiUOc6qURztp6z8/j+J8ziI7Y
j40ALc8LHhv68DlZfMXBKq18sSqrg9uYtqUyiD4TD1oMtToRzXLijpDzXP7BfyE5jVWIrOThLt2y
Aqj1OxJBiHTeACxQ/R5xjsk0v8NIow2P4+tmxP7hlISTdGDZvQZcLVHc/jo99fKZOLQY9fJG3izE
SkZ8VvXg+iZFuYsgIHX804ymLP8GrkeOOg4tqXxN2jubAlDGeMnYDvFC9mripmOEai+7oGRwVWOk
FAxHfVhSn4/5imV8QhXUG0M4vj+s1x4nNZVIX9fsFqZwRc00rxEO8KcHQUAZtWMr5fE+CdCXdWuQ
8DROJieH/LsZZMYacqZ3kF9LyRRS0JE7x8hEuRF+w4JyqvEq4K4CfpuFm5K0A+pYekg05LqLjAHG
o+FQBchubp0yC0zKPEmMGLGbN7G4+GJvAhJx7n9dtUEIRJTya+5ig0ymNeBdc/w5tnmzG893smeM
umH3k1OWDNZ5q6mhfCQdxOAaO8LiFA9sgXxxottG6VmvkYi4pEowUXIX7EZJbwoj+KhBx4yeVkPj
9NZfcaML1UuGc/TDgcpdcfs3c4udCVrQl8JJe8KU4VQUb00qhbz+khg9ghydNwOczWwHC+oLzLya
mUsuzXGD50JfSN8rJQPUxMXgD3/f+qkQ+RCvSxYPF/Y+gnV9LD7rsyGWeLuLeqdukyLzZ3i6CsMy
wfV0NNDJh/dEVPYddnQZpZCg0XIe7f1Ub0Bg8sG1tQgj4IK8XxHO8dIdPhxRF/DLgUSMziqQ9eft
GJRHQ6/PwId0IiDiioWV2jsjMFYu7I/o67ODLGlyXAsGhFF/Ch+litg5txDJSvdxXSVAmzC91zII
SA0AhqTBop/p3sYevrLJm5Ae1dhf3ni6t+uJjwIV8sMujY6Bd3hfg0xirKCfo/hYJiBU++7kbxt5
fP5sYVfCmK4KHazwE4P+t7JAPxffaFbwtBmS869GEaR7BZ+9VVPT+0+5Pa9u4+exVA3i8ErqizZI
zXKxNuXFr77ZVD1k0Q0xYB/u4BvGAzRTEhVjhoBZLzvFFZQpY063oiTOcDaO11FqHrivEUGsx0dq
dDgPhtV1tQOLVfnS5sowLPW7yj3ke+sk5UQEfO0H7lgNveCkGTzwYA2FkYPK6l9mNHf6+ppGe5c4
ldddXMRB+ClJbvftinahXAodtH/jkK9Eyn7fWTvwS21s7LV1UtnCUyEyngivzvcxZfZPkwCmCdik
Wnv+Ql+G4UKWn5wc4yS0+aZB2nHyZPUqO+CE4vMHan1pYF/SJ5QgIiqyE5lR5GdXEQKJL41wo5Lu
hvFQqZRArMUKRTA2xABRKV+RR//SBnxcSl1ZdYuG2i2tViPYr68zEzeSi72JSTwf19DgQxA3RsV2
Y3rzwkQhGYlZL+bC9ofsAa2VG0uq065gy8u/U3nBFVa/15IccyxRLDm6uCcKFUoYqU4AptwWAxIQ
U4DhNuQA/J0f5LjVO3FQ4jYJtNgBKBt+1Pw4iNta+3iANohw/mcqn2SNZB+001OdWfnDP/ys0OAd
LsBHfZVUvIaD1GywgKrFDh07EYt4/1bqeicMJmv5PLC7nWgAFoqzkTRRqFx2sCIf1W6xmKPvlDN2
QLDiQJhuzyWnp5tekxFHnO8Lf99PlqiO1aQ+qMkCI9ATzQdgYAk58MsJ9KoSh7INVYOpJE/NGe8R
h3FnxkIflnjYh0+wFLQ5J170N0yuIa5LoadSUyEG47dGwYgLSUWkiGFLX68K/1zDs854sttxS6Ke
y4saRREUnpDmbF9agmcb2kxGhhWfctTI4lUJlqbhQvCKUYFXx3c6wv48P/HQPI5zkLqFWLAFVGpU
sUG0I4K39mUtxEnA91BEk5oMf7Zvm3/rGPT4Vh5waYlS8WkL2pMXtWIokzvIPKEi8tVK1Ez1wTfO
RJB8h2kd/myQf98hqJS9xkmNi1vApRzIi2VH80G/WWWc6NKDTOGzmrdi1ssZGqabCAYOwvuifP9n
hI8NSJCKTyGdrE+s2WxwWTAf+Qbjm9Woa3l+/wpmoCFihDbtgTttIVVLJLSpVSWnH9p7hlGyaG2l
C4Opa0+pH9CoHKA4vc01ed6mQnDIz0ep2MB5Gw67x3lCmp6ViW9rupDUwg4opaby4quwNsJZy03l
GIHEJ2E5ABoqt01hLY/AfwvqWMaXOprvnF5nruP+FUh+VhMAwsRsWDYzhMGrEPZhDQYe0aWIg6Qz
WlXBdZvhTfoEgtsEMoXjr59C/XvfEqlusJQCpCO+dz4qFt96EYFQM07m593Z/G5FNni9CiMbQW+4
jWSU+jXKQRFwXHdljKEUP/kRJj6bHV7j8/t2HR2LJgeq8rjw3YBcS058ckMHlGtug+ERhda+BVGh
VCU6vvSRl4rrDw0iXoC0a2X1YqUG46xRSKDWS2HrC67R2oTVy2Zu8UNAYvxdUFZRsqEkx0pwKShp
wsWAWg2UvvlVyXSedt085wn5OzM4BaMxNyVSBPxMIzKiSaAVJVpGR1TTQKB3NEHsI2S7IbFk0pKN
2e0m1FSTjpcII9wfxNqqvUT4OkZmHnkXK7XKKldmdt+QC42hYfVDUHBvqdEDAZJ9R9/p6kwqwZIR
Bp/o2AyxwK4ww+5oNVNRHAPxfCOcKbowZqy9/sB0j4/tIvq8B3KvcC19sz9BPH/Sp/beX860c1Qy
jJ/IKfputN9wlcbu3s+Wny0q9/9tgAaG4sFZWvHEEVgnPDLuV1hipJZ+rxDfvvmaI+13VpDeOtFb
qC+hYfICKVJFoA7sx+2LtaJnrofdegrXvynZd//r0ep6KHurZQri3SElo7lzaRWHtUENwvynHrVO
9vjq9IhwVIh4oxcrNwvPAJInjf2LrRcxrohFM2Pg4qf/ZMDn1gnzjU1kaAxr5YKl6hnCY+XYhECw
WMJUNp7Fab35cBo+da/HxDQnlcABAgEgLemd0B879Kb/+e12fQlHHshevX4kh0klgBVO5ECbSTO/
EwwXjPu5H5B+wp5//Td1bm8n8MWXmE/IKXuq80CGHh0QafNIONGKJmts9qT230/8sJFkdEtC+546
v7JV1SVvhmCeoet7k2KALXEKasGjCGkhMXi6Qx9HTtY6i2WeEfvdAk9hqZKPLYzsHN7Xrp5bwl9P
vkiH6WYzrkrR5/HG+tcK86NHS7eJt72Ph4qY5sVZSz6Uh0su+3ejoxLlsoOqa4BZk4il6fOd3QsY
0PEZOLI/P+0wmrcvFI11hxV/c6virERy9TtDPig08H6YXh2FwGgNCmFIk/YqnywT2gLWxER3/j++
5Yco0DbKixfTH04lr44oRVoODp5cjE6ohWWVfEsWYSI+bGw9yb3g+tCFP+hKbKZeekH0A/nLKg7E
On6Mk30ZKXlT4LY5ns38nhCRRw7QXhrDGDdlcY9gpf7AWqD3kJGYcSvciM83u4yvbSFOp5TQxKEc
LUGcv7oznWV/wQteWK1amRT6VW9sDpY0MUZVjyN/wwWPQWaM9XXxjkPHSPRe+GhX6d5AeVpkiUzL
iW/Dv/ES+yUap181ZAKJYaQUYWjsKiwRXPq4F6RfAVyGkhGGRXC7Tu91bqu2C/HuFL5gUIUP2t06
JlmR4/3eW1AguQYRGZX2SWrjsxDd5LTqVJ1u9pEHxd4+LE6dYHHEfb9DTj/FlnORFpXZsFclqZiU
UyqrJUTy8PUxTU8NCb1uOHIKwWerClRWH+RDcjiStkEXwJxIEm2RKeoPGv38/VaqGLcwYi7dugBt
1Q+etLqLbKLr7IlH6gIV0nZ6bCLvTNi+WN5y0U7d8CAMtEchzo5CrKxTYb6dQeH2DbPv5sfEVntq
6/KkpwrrrY+Mc4hfLNISq5mOFR8tzi/0k/O+gAdUZLEsMJ58nfFB5CdQSYYaCIhLBn3G8wMlm5bB
cJob+nwsrotbmzFvH9o1by4uGVroV8vcCkN81fO9sV7kHFRW592u/tsqLBBSdqVYm8QRkWdbvunW
am7CrdYkVUA02MOgD2y8TxhGDCqXH/zrPJZD43LRmGlFhhqnsaCEiAokUIgaq1bU+sGRhAN03gUP
lhHEwTVFo5IciWILRtHh0WfboibafM9y+W9hZMGsrv9jKhL+Fs+sMlBDnqioBLnGy5IhJ3UP9Ni1
mvHPgONW70AQ/bH/OQSUTrfl5Ra4vrJKEcMzwk/h7xXhQX2pzSjWQQIfZ/ZsRFxptEHOltCRVp0g
OV5/aYGAJK+MUD/wsCWO0nxNAuWyNaeE6sEZqKjGu+MRP4elE/R2rPV7ByWTlqMWKFQ0CheBox31
iXmPGm0DMbBtnn2p7+fYEMGKGZqQcKYYsItsDmEkPfMn16I74hdSJT/QCD0+qD6jrq7rD9DuKN7E
eoZcNqKlje/Jpk/0AQJWTg9AmlvCqVd7iornQYUysHGvWhN7A8kT82Tz/OFsiKJx70zQNI820Wly
nVYy5MMW3iDNFHU7TVl2FxU3qiMgwFZWtK2S5V7g708rfcvuo0cjwMPz4YECQ9zDKz8d/AhtSqbu
Z0kF0dsT/iib0saOpJ6G126dmlXVi5U4y3Iv5HBGjiSDgpIZMnmtGtCo/fe8sKq+HEf+7CVRtFqe
xzfrnxU3Vq4Xak0g24/0yMhznD7cvKnpb8X6HGNo5vX8/VSWufF/hffYujBc62z4U3WgMScnJypR
dggYwKDJSjR9NgE3BbaJYWUMCI7iJvUwSnbOBbePhTgXIEGwyW5ABbuTe0/nyzdfIiwyopW5k2jm
4ZhExRLFk2j6XVNvK1O9GXLiaLrChjE5AnwQqtZGLbktM1yGb+9f4gdJuT2/3vd8qfu6G36hWqI8
hm+ZldlfTPlceFkFizpfOZOj7q2tyYWx5x46yC9681qhOFQywQeU3+h+xoDZdKDY3Wm2ICvTA3h/
nrk5mBoRTtMzoy7a2xG0qwL9UadpQFMniCvBSYiF9RhqsxarJcW7+rALesoBRkfvuFf031FGXLDB
SoxuSPPRONWQGLkk6XJR8iUjgQHVApVLosU8Z2WhDL5r5m1D/E+LgsJS42ADOhihGiFjLbb/C/Fj
wkR3omhq7B+v4w6/OnHSS2czWF0KIKd22+5yvrIy5I7CEWVKzssJKVS3Z2MsitB2K2SWMFCWCGwA
u7NkcvNpyuMCOPrz2mgN7GuLybb2LWP5SKVlVR6JlMQckjq4ttrtXi3wwld94d7RjVBr/blCC8Y4
ZJOQu2Hl6PdgUPvdGB23dhxc7nof6bMTdOBrQsEpLOG+NkVM6631KWuiNG1JcwKCsw8FnuFoGMMN
JHrIiZSFpn0cU5uoRS6Psq6wAYXMQXxi91xlnWW4KvUW801fKZTzqlQiAmjIJvWKGhc/rAITwjhp
IWVKfAP0xU+Phz2nFeRm2zNddPaZHhwdAkBJmVoGzH4tgLJXoSp2KEWilNZ0h8iFRrKMbykbp6EX
6krblAQoxqipMD6ob9N75348aSy9d4931DLf7PmVe5etk/erruTCklTz1vUu5pkpExRdZHjaE8YN
21NZ/i7tYByHVT+oZk+SMMsr2rwu+a1pzIfkF+/vmzIYFjYoW6I28tW7MXNpxgoJPcxe5tl8SSWR
BS1xhAbxmsHl3G2inxc5tpZ4St48RAB8y2adLZo3trawOu8PK29HXX6kO+zVavN9eqB7w/D4kw3u
r2fnSuFeIGivBhbhPAUS2EOZ84WyzukUz82d7pWBcAQStGajcXtJ5jYgGyOJQYJ1s5/eDzMe/VZM
uxvkB2OPxV2k44AxDjQ7pFgr5GG5YZFg08fE+jAZMzN+j5e1e0UrvsqXHqbPMEuypHUtBUEVYSSR
9C+Krcy3TUfjO5WoiYbE77Y8xRBJ9lSMAvv1ZFCt8Jqh3UrY+kECo4oodC2upeWN15hybssws526
mKwU77rndFAko+8XnGCZRSifP208Ts5Enlc7f5FvQ175H+yLAmTy8BDq3KGgp8WHRVsEvR8aOQIJ
EiLKlqNZLviGnd5Bxh5q3aDTceHPn+9fcR8WHxQ7MHlmJv8OfewEwbvgLvP6ac5agt7E9LX+zR/W
12OjaZ3E5/Hrgk/cqgbnQdXkdektNuwKY52DebP09jzwNnXgdHUdY1UZRwz/JDRTyVbyS6mkhrJk
WpL/lj5KStNoWr5jblsemSl12v+grm8a2SliZBHr9lfyJgLWRnyR9GRqU9SdsI2tJShVEpRuaqB9
LLqAdBdGFAFLd/pC++PasOM+CUSdpeBqlj/MuqIw7Gjyc3ZtrHfv6o1L6TpVFO49/IhFp9SYpCN5
ATtPskG8MuFdmmr6S26yWms/GNAb9nQEtr5V1e68AqVtPO47N+jzgJP9TUmWnEoLFIoSn9CWz323
mt+nh8hQsETKnt6al58ETvQg57j5kX/fy0H+A8XvIqv0c/PJ8kVsG7G+4Cfn34rYEALFTuOmNaTd
JBndBp0TSBxLPLabwe1mQQ3IFKrjnfFiVDtvsPJRZVji7WuZUeCJTb5bzJzsKUUe11GL0IrOwwT5
CdbzBxqaTTcotG/URDZjPSnQdZSZMlGUkh0+EQSK1chB6xwYzpaRImWYffhsI5f0b2bqhjxRt/Nf
RoU4VmN2eq39ugUZrzVuzQc1MCYgY1CxEXavG8DHb/GFsfkzQmOK/OzcjBhTa+U9aOw3Z2y+Pg++
4cT7TSAld6BqQHltDKMaSTOBs8fnq98lSB4PFwfvI3JsQxDmsW5O1Fp4U8Fp407BzCtFU6Ru/6zx
aWFPe8gBsrI6O9TlCqfnNhGKeP0yWpr1kQLhgQoRQpX1oLQ8g0qQDHyuuEnYM/Eckz+Euy8xMlNb
2KhxT6+TrD2eoxjh6k07HMDEZ+oBnQ+fwZ3HvJJKn7THa+YdFGSsRYqYYPEXSvqeR9GVGCEIj04b
GPIedPO6yDW577HpupTCTLgcAvic0G8nAASXLlXODNG/Q40Zpg8I3+9DmXkwfYMOIOhSw0iNIbsN
VWMbIRoucf9k6Wh59i48Isj8ijYelP9tNO8ux/MAOxSZING/9zkOki5iubp6tn5kW2pMn8t7BGN+
2Hagq0pm3JJmlzj9Vpmcs39bbNHVhXHXMsr7H3n1KkSswgbuMy9V/acFYX9ER2oo9l4lh5mW9P4+
nDK0O82ygzgwbdksQGjo3MCBk3IlnpDLiOLmXNRiv1vtbj2B+3mHMBWcGn2gtqKwLMgptEyxLdxz
ohz56Y+PRT2wiWSvroBaThtCJ6Iij9uHzBxNHtlvPAgUT+yC7wU0pKl9c4oRuwolTxf3XwEnrlZf
kz1HeFq0dVp0o11JnGF7e2i+dDTZu2+ywycBCK/3lsVzvmilz4pQFv5T+avP6ASe8uH8DLzKTEIK
hTJDNcYgYdVy5xYhRvWii+gjwpvNJlS7xewfXcgMxdFPwrYMc/bgZYPx+1ApeEdTN6vp2lKDMl55
43k5ReYR+DNB+eXWtm4TdZ53GNQSIhldsrBVpOgH3MyTtvqEaYyMk1T2LJEHWBxQwngzdRlQmZCI
xds3lUWrKKFE46DvCrgax+MqkBlCPUtfI6zfTXQsvs9k//mWQzpHTqStHHCJ1NoVPfNj2Tphyiv4
L1iiMYNjugEwgxO7iKPtD/GisfTfgSRr+ewMP9sm+Iq6u5KYCz9NiUycTUNRdAYXXR2tNlAOG7Iz
3/SdrsZJYfnpCaNMkMhJSZB/5vwCJFDuNVT67uLr/98Bxos2+Gv2c1sAwXeIh/ShPyCtwC9QsF/b
FxtQVJF32q9o8NOAY/6DmPZ51xY512sCi+PTnhe9R9kBgqGYpfV43nLnTgLoXMlVJkOEcuH6yGC6
lC2lcWk0qIqpbEHQLJeunb2VvgUUpOI/V5MvCXY3Fq4YwjbVeP1v9Sa3o+IHoAogCeez1mV7T51Z
UY6GKcKiL9K7OjZCJ2AkGR4kzv4wK7YCW7fbNf+wVWskua+r1zP0YxOqAOzb82Q9srAWAP64ePWf
n1XtAR4PgWVfiEgCRAWwTJ2az5ydad4rHHv9AmwelscdSqa1MhOEDzB9q577+Xma+wA3GtvAcDCD
KWOoZot5DtfeUlLW8MBU96dAQ2U4lkselld4mDfrGFKc8jAVJijDLqEVECSO0QxTO3okXEHZzGik
8ZeIIvbdpE+C/zZp5sdBK3CkfKtu/qI8lPdVd4J5i2bZPDqSmQL8ODWTdCSlXG/Cmm1KwMMUCHKE
OyMd7XTAawKvDzrOL6hk6djQKQPlrc1SgZh3pzYpa47R+szisOCSzDGlRKe6Een/N4lExIUj/8ow
N1aL5EV7npJOw//D0atc0nIS9Azhuy9TI1RaKxjzdGXj3kvEo87+yWEaDjZIVoLlgbleRchHpai1
usew9WUQ+vgJ5zTW77Jr788KE/iqBR37UBRJrUJ7mMv19Mx7nIMt8OGypvCs7wvckiOaFFD2IBv9
YvDvmqt2ei890HXPCsAR7xfDDoJd5JXbSAPihdlBA5Sk6q9b+zpFgjQz9zEMyD9NfRamRubQi3b+
UMuVH/qvEHl2EevTKWLuGejY+uvFNZ11saWYLFgSLgMiexcA7fEnkeQWMJCBwEnqS3/epEVPYUg2
xzT+mzJLsmHL7Uk2wLSH6bc+sanqaxfJu0n7pkSaKRt/fIA+2ZuKpupiOaR2j6cFoid5x8Xr+5Jp
adSC3akZepAc0euiTW6SxeW5bPYP7Px9q1HH6HmO3Zgll6S1R75mLvAi7H73eoMfz4N5GsuW/vHx
8Dbvl3zsCeKr/OVKTLr2cjlS6Ge9gHOewHfZoj1B8gnocUa+82P7BeT8AhSXPX06Wn0Q2jJfhowp
kWPEjcHrlvU2nNtI1l8g1/gsAUkXbb6euK7FMq9ul1n9xDVECgTqjpUzSm1GKrbZ91HkOf19oP7B
0gD/KTPluy9fZKuWtiEQ3UYXuTBpGYdtxsY5NZD8LlHSsURO1e/7+FdRTBsKAtOY5JzsKv8JaEvv
Gf77pF0J7tl77nQRXgnvqeB0lb9u3/oFrAachmpdWSUiblHaIoZPju0RGLRTfqMw3Y1Hag66Se0O
1hdjF+gKYYM3USyiCfQU7zZtbXu1OQDg/LhAZVPlVqMjyp7SptxoqIzwVH4gOkWP0XDPv787Fi95
nAHT+eMWblSZly4osq1vib41KmM5EMsTo6j0/BKGrSWJKLrSerLBri8fzpR2djSd6Z98gArmjsCy
45ggnGRlDLIUnJ39KNYliUWx056221kXJ4bfsLuY3uLOpPC/TQcUQ3DlNMmaAq1HTVknN5kWlAzD
Nh4weaIlyt3AuOI/p5UtJVS0RFPshPRrvHniv7lzpXKD8pmxcoVC9Tock2KL3pQ1G4z77u2Yv21N
JLTMjB8WhJtQfBznQmG8xPqBPuCoqnLYAsxpJMPFDfPlRj5zY/WK+PjjmKVGtLQ2dgPcUiwSS1dD
Z1hOocwKgSYEZhk+38gOzz/8VJ+7/cXMSo8DmKgWPsxdlYTF5TNNv7W3rAqkIeUuENUPd5Ai1uGo
5IGpj8AgXjWrmD1nKwhZSgyDtU+NK6Rhe624tTxng/cmm7aLRjikaARpkqA4H7e9rND2nPlQV5P8
osOfvDZqaEM1a9LnMlVnpEzdE60kKBlkO3FJuvIAyDq9e000o77Q9wcvh5JKpNYFUg1NiFA8n5G+
H45Pb70k/UT0PlvZBSPtQSdSIGLZNEjtBOlQvAFFIa2ta2IRhNYKbd85jRRNLOYCl4DtFFBP7dwY
b0csv95PfzHEqe7Z4rTXUXuzNn5x7vQ123biC7yk5Avy/fEt4XSVYt9vhDGf964B7hhNCkw6qS9o
AWLi3uRVox/IzcWItYTNiOCdZwdWf08oYsjI0zHAplWQRL60M0wZGOj9h8vcVEWlBnJsth7WOvWT
zSXEI3GTRVDleV8xS34MLM4suRCaU3fNcoFJzhZUoFh12wqir4J848YFOqVwRVOYMQ3Hk5AzwFNy
3Wjm+VFJwPOxNyzPZUl8wW8vZ1BWe7ltIetysqz2Nn5TCsvJcSRxqrkoccpC8SInqEXKGzOeHVYw
gXwOf+u1GqpGJzBunOpZ/+FxRe4sMTxcqeI37x8roY1O1HHhv9wMzpV/zH6B/6q2tQI6xjWOMrp7
hubrUzeE9v0g8/FnJxtom6NxHxDENlGdSfB9MhDkdNlTslGF4aMcmClBrgMlBZ3qxyrOLMIE7eIb
1ToEBnJ9NS9OdeyjlLbaTVTW6a6QjaOGtXI8Mh1P46yxfHYi6igF9fyOGlvBEjEHWWGTjxxe25vL
t1D+3cETpuaSAik8CT6flGqN79GvDF7IS+6V0mFiqJSFEiR2kack2U2gd6wjko3hgqbJXYj1N/sc
6WMuFS5sPnrgzr/9Vzt49l+thNdwWlknvg8kwzs6ReymlVsFG4sJEdzfqU0BuN3DLkAfAeNkUmIz
lxnV6hdmuNkmzlX3OMx9SzicAkhGyyjzpIBrlT66iXM9/2UPepdUjD/yHUz1MVZe3PINuqmKa30y
mLMDKHpHO4wl0+ni8LPyO1FNNa1prxhLAj5wf9uylScaFRzHBwxWN9hdIiTKv1VBvFwbOC836RKq
nwYFpihePna3O7Eoov7UhgOq1fmC5Q/UoUYRchEdLeuRQMoJwPMicCk/3fwvuAocqLgy0bvAKDsb
OP0Da2ay+JFZY5gdlriT9CMWpem+edf3Z49/AzXd9c+I9XRXvi7JOr7leritwK89uXgsm03NoJ7m
T7jOPcQSPKScZVa8/GEgUm5kjFeQM5t3ANycnaiUgoCDdhlxFYZVeFjb5XR6UBYoSAt+FS76gB7P
vISoNhn3zAicH2gd0VdhLQINPcD9A3iLLhdx5yZWExGTR41Pg3Uir97sog1Yl+SyCeH3Ire1zaZ2
QHWaUEGNV7kYjUTKxz6iB5xVdE3xiqvaFqhPYSHZAD2rur1fLVCCNwm/0Sh8K/Roph1Cpnc3QkAR
4RMqh6B12GfFyCQmpYzz31XMsYuJUejg5mvkj3P3Xd7arLKnY9l49kEXmxD/0A3FYkw9fKrjqXpC
GpmtbKVXp1bvH11ixIb9oCI08qZtb89npHuEe6rmfVfElw+KlPB94aAA846pW/a6vMWscRLDEVF8
WZDljwXVF6H4WPM1i4WLavNppANXI4erNE1BSRsLULrWcRrV5y79/X3qAieOSZ1OlFuYM2FLKJb4
G40cVlrxdp86NaVxjZPctndha7NiiR0HXqf3BHZsA/7/+4a95MdRUSf8qmAufOwp09aN+0L42oae
UpnYT0+E//LivU+l5Yi7qbIV70GsprccDUDL/zj1E3lp5QWSjoqfXg7q0k76/F4qebi8hXh0N45g
fzF3U+0mfduB4Y3B3tbJ96SK+m3Kg4ZNwdFuxzsDTzrchW2nL0wFpzxWB1XkBBD6dnG9p/HkJ2Td
c1H6dloE3yST5Nqwz3UNOkyCzBFiuOgMPgVI8L4IadNw7tIBcGrQZsWZplknrrVixIcXYfJO5mpi
X0Ec7LEBHTgl50CbnPbt3NgG70jTmO04IrObH8OCrdTCTvmY5SHUVEnkg4Hc3GmjDvVxmXnI/WMk
t2BV6mlkobU0kh0gwTbQ8Cen+jCtk3bN8HrGqHqAJYc76fPmYLwL2ggK+GHfmX0syutyuyqlJJcy
ss0jembkIea81kTC8Jn869UKuq9QF/PklyEkVjV0sV2Pc4FoADO/6eA848pY/ndeyF1+MFCIGORb
GMDbeYH1b3yCefp3D21Dc2RTbiO6pnPSZSt+dUJKohWRH7av8Wp54w2+/rZ75NuQ3l2XtiFLag0Q
F6FooTacTPRJvqDzuGEKcPfGd03RsyEBh97TPacR1v3PL5xxKeQbryObxdJ9VH3pvKIRDJpVInV1
W5Wgx4HrXyCKRM0w8RKLut6OeIbhH/chacd7atZn3HD+AbN39CfyqDT+WMs/GipTRDz1j/8K5Z5f
uBJWCcvn3LEMiyVjsq364U+SRdn+gfsiqiFAPu1u5bMCdv9gUqY2zsHs15wOkcb1BmRxp1ILs4og
h7hEdDVPKyKaUaAFaId6somoFqMtI94kdW9yUpxTfngbXCBPOGWdXx7dhHNUATHbCYGnt7lUeug1
VjIytmLbBLSB70EAWKlph14bbLHcAO3Or11HkmuuS2Wx+p8569UfGxnPHiPciL6PlHZwAG3rtY9z
N8PTCo9Prfbu8FKijICSZQYPNTxebb/eNrSQIk7ImYnuyOFGu5iMoz37LSTsF1Z2lC4vkcVEGfws
JTvt95ka70qoXVdlS2JIBTMo9/MYL6ktC5UFcq4ad1f6I/gYLUGlsKX6C+yg7MqXYjnWPuRKtUcU
1VU9deA1fc4x+v0tqJEGxKlmLpG+W4Q+q4GQW1nZ+Ny9ZFP+qC/LMXYvbeHwqnn+nOr3yp4EXQrO
K54hvHzFvwuoS9TnAeBIJJy2NyHKFToYZjh6qQZP0f/Tq9s6rV9YDUEftX9n1WFdAOcQ+LQeVcN/
+nKunLnA1ZNC3Udi02vdW3BXKdcCsgTDiRBxNRjrcyxYlox3A78SpqLDKPsU8Ioa2o+/qMs5TnpV
909Pe5K/ShKXZrFAkkkAJtfE7MW7CujOgaYrcdja3jGEJB2OCUwmTtXBnfQrQcEiDbY3uXvIxosK
r19mZ+XswrnqjcUyaLnzqqFtBHp1QgidihXILafDYCGBb6ykBbKSh1acyzeCO6WCN4athd7RmM57
u/MDkp/QZwWrZ4xbzx8QuxYokeAUTEd0UR24pFaxWD3KPxZQy8cf4banW+ywSzbTvCuX3Rb+rz4r
zEWRAg3h8qzf4LYTmTvVkzAF+sh0fApJf4npuhBhYMHeKlCgqqyOdZDI5zzZyzsCooartWPRAywW
wr6q+RWM29B0tI4BQ+jpsCz3zv/A8YQep5V/lVfPYtJomWJvBZezjH2uvBimU+tlhMrlaoYd+VHd
xlWTbhMdd91IIXVWAOO2S7nsQKVI+qBmljppCisBA3w8M734XBXJzegnJ44tBHtd067yeO4UFIyB
2lSPMs0vIgpZ4qR8tLovfkSjxeHTcjIumxhFpy9ErtIsnHMWTCTJ5eXX5wWmMq8lUMMX7Q5MDGnV
RBruIK3f74v2tCd7+a4H8rA3ydAxlc0z4HZkmTd/xfe7WWsZw/RKqCZVLRqhJXQRYHDZPcYiqC7m
wmufs0w9ewPw8e16UBZRRn5TSGWs5koF/clcz8J27H95DVzeAO1CXdV6H4Nvp+ZQSABRuCfZpah/
RzF76KfzyraM45hsHyHsI2RWFf7kczpY3rux+r4W2U1PcFAc2qqN6t5qsLxPcBosTwgz1JiM6uq6
qMvaLyF/dGqSVNQFCSURXSfxMHpRQigaQPEM6GMbCFE2qIof70/DvkX8fqtLSKB9TV768v8YtShN
uUv8SNdhrEXFLQaPpzNR5txEwe8/0wb64KI7/dptERR848KFth+YzK2xnp7Fvl+iIKYYQxR0WYk3
3IY9lhm/H2otaZmsN7qE5UGE4UoaPFBR0aO2CnDKnDF4UGCjeJSAurrI0MA51EptMb5DoTJwhera
gCcM9HnWX7HNlhsfF5dbWKhSxC82xA/GFdR0VFSMF1Z/VKFD/DlIUQOMUFZTkY+N5WHnw6Epr3hJ
LepcyIxWNgApZ/ykGNa62rEwrOHVxTz35aWl1bHctrwnAqRO7AKGu40rCsYXNnpjbdKG9LE+NkjA
xfQBjF5wpbH4KciZPtOjGcc+jWR37/sHtDGLjCrCZN8A+yEUpNSk+axq5sdDyHESrxCIjcPZ+KML
zmtzgxnc3IKkT2OLkoUwFZAUCBUykChQCXOo0xezigffGThN/cYFvFx/y+oP33unfoYawlqFigN3
hFLGZ/tBh9jpU+7GiLxEp0qkWpTnJNehfK9Oh5txqlrCxGWNQBBXRao3jgPoTk9D23j9T2s2AX6/
giwz5S4h2TuvXs8YnnibvxWbLTQLeLCZPgusA52ZoMkC5XD2KPrM0sRx3aLLgkwXNrlmB0yGT4QY
FM1Br33j76/+F2qRL26Y2oftyt2fA9MS9wutlCWMkqkzWBav/famPu92gCFaiN3Ne0JqvR2IhzIo
dVnOXfupOIN/IxEvt/gITseeG3Q13cx5ZaFHmsdNbzbmv9dw+v/7PTDcvudlfRmSa0PeNfPoT3L/
xvyG5jQBFcpyFj/0C0tjpe1hYbC4yN2V7w2qyxkHa4MUP6KEHedByySSwvR+yD/0pGiJGYqmQao4
cdEUNUoIHw19AoO7+q1s1oMFJVnE4hvqcUYfg8QMPGlkccc14lWKX78xhLb6n/5vsmcJwnDd6gQU
toopece721abMAODqoGmgwD2Ng8BN0HvfoBaIOP/ednfziELOEOpCWM7kFW233CEf+HKhqtAzKD4
EPt8ixF0seU1SW2nbBst3nRQVpzd1odg/vq02F5S8fDoh1HELNIjzjh9r3BNUCQxWp8/bw4OMLqp
4ce0+FR/5L2BdDTRgZ/ZFcGfPeS1wLBm/2mDjX4q/CG4NmtrDPJ+qKvZqov7+WnwCZUSX6qQc41s
+iiLHwp1HozET/zbM7CWI06BinEWReLEdRyMQOpyNxejWKDkVAKWLr+NIBcn7B9J1uXTFpG6pzp0
YZG6HRSO/sVxbH/BN7091hxNvKFW8fZ288SipKaIspn9VCMMZajDdyPKxDy4ucQQj0tVY2jY4fty
jmvkJIHbN3cUA/G85O5wV9q9dkWL9n5v4/nhaN3aIoQJFTSCuNswvF6g+e7/ycWZlq50zbEaaONb
CMbimHD/2pYExT1Th83hHEZeRoBVwx4RID7lxHilI1xHdPIIw4Q+UHz+g1ldmuru2wJZf0Rf7VM6
3OTIZvXuGoKgQCD19EezGR6Xvz4BgBdNf0M2r7lm6MtB3a/NDipNIzgLOccZOarPiA1fJD86BHMb
6q6OWoOTPC1fs1u9auXQYtBqdVjbBkGc56EDnlg1mCLh2ustt/4Fqk68A89TFMnq37bN3vmlEjav
6cJIlaV0wu/FU6Jw/CJ4KX16S44ju8idkgw/Xotwg68ikUPNBREv7m8Pa2xVWtonFNwwhjTyqxde
E5N+gOosUGHpD8sChT8/BaV6NCI6bTWeQMLPNn1XrJm3LvNyqDAtVtBMM+eeRHLhpe3AO+Qb7lqy
c/D9/jdW4mfMOwp1NoE5VT4TVp7doeFowiTmynyoOqFFgnIrH4DAjk3hmUg0ePBQil7/orD4u3o2
T2KzJEex5X0dB/gmvCytW1XFKaGZe33cyviA1B4JM1MUQP+EFwpOh6zf8ibS9XFL1jVKKbrL10Yw
Gk1yeO+S8asBtNnqTXH2HfpPZqk3rqxAoNQphTY/9qn4Rxf/khz+1myyU3kw3mSxBPuVvxURW/wV
t707Gj7R/IkGW6VxRuXp2kSdfQR6qFKsFCxqqmkaMtYimhblz3JCkE7TtP3hNL8Y3bxBVcLJlxyT
AlW0TOEXgIQii97wVjwG5Tj829lrra/PsL7+nxGM6fPpIMiNoIZoZzMNgI1/9CCWYMbE6Pdl+3Gh
mzsCkjwU2w2FBwZoE8wPxL872XxPV6ewZk5Nztz3oxUUNPk5GiUadKVChC3qE4c9WBuxnobtzkEY
hcDaoK1xLuhLq15Y85TC/Q21PhjRnBcFQsgBgn1HCZdvYx+HNmfbYPt0HqxMqJH5LDBKDPM/hmyx
OoH2OVPa81M2FAArsnruPoGAWDAuNb4o2L/iPpF1n2rGXXaOCon/rJyB0rm1Rg38uNGd5vECuzxP
N1gvJN684dWhx2fEkY1HrUHxkiPrbkIuJHmVV1Dg09F8NmLqcEiXi6e+DvbKEYZb89srI6DRFyqY
CVAXVzgobVShwKAI8JviqGfmHqop3UujKFcK8CT1zM5qvYK72WfTNZ/5BQjBxa3wCNycXijf4OnW
fAH2vQAzmyeUZ06X63uiAYnxF7eIFYbWFuHr4KRpsiKek81W3BBjXT0+7aXBB7OaLsf6S+CHFT+K
6rqtrChC22F0nXQTgHqCWrhWaA9W16wnQHXMAIPnRKIKXYniOqdgyHXMZ/8LQKYK9FOpgxUQ96rQ
9FvcVy+64XYPp2OKmzzZwlHBSqmYpL7hB/clioXN/1IJRJeX0iCe4zSGzE4toJynLUYyDJKqPqWb
Lnhi8eaNA2o5M/ca19w3wLAwbuPvtrAnYQ5DIokDGxGs/VUxhh9nIkFgc+kABKDIIc8oQt+wZKNX
4pQzoer4RuKo3cen1Ot3P5JTwwsyLVDzMVAjCXglznqN10yCCK7L7UDG7tMOS46+kdyiuY/S6KwQ
hi4oFBzESS1TeqrOUwN9kx1d6mpaq++WM8FcIHTq9gyWaxszWBR/W7zIIOdyCR3MuXNlhl6EVdoZ
6ROQteyIIG052qOGtqsbh45Iwo6QAToLbQjw4lQHio549KN/JDL+B89rReDCGVNkF84dbnWo+cPl
/oWlHGt2rX3PWT1LHhBWnlzexfnnxDzUOvNAA2337T7lLuY11Q63W/Vjhe5hkgPjfTXLDomyLdMH
JKk6gYk2tyLiUG9G3QrLqDb4N4sYgq1LrACXCbNMAbsl8Xpsas2JQEO2AtVJPbaLGKWeOADlvftS
r1we8bTGj3ZWAthqTDctnbMHpx+K5UVj4xwvoSr75FaKJ2yPKhxY+a42SgQl+8Bw3VRRCJnFuNtE
Yer9JvNehtK/kMnBzDAd2UDTU6FAgoKg0Rpk+ucsVOJBoxhHristWwQVeczlVKun+NYOSAYyRQkY
jVwuYjPap5yHOWvZopN4QMuAKIAGlVBeAJnkvHt7fx/7uEy0Dgi9j+0TLI+9N/ZEe28hq0ykEUCX
wz/49D3ODeiDSZd/9RSb/sx+HLlZ6U3UqBz+EpsGAG4ASd3Ak+qsNivKIflD1Ru7TsqEsnFTWhDz
sma3YgGtqVVBldaNGwW8mbQxuOKnaVRDKE3Gfqy6247lhAzUMj4iMi4uOueyFj/7MGxck+If6WdN
x+46JWOBZXgsk1gqvtdSGLtttllsI8L8Ae5ZHVOr2oW3DKSFSdQxmtPDTJJ7tBPCBDxoDel1CGed
Ly8m0WNspas06p/XhCbjsZXFhMikde2l2/3q3voVotZ1C7IPKJGhvirF83j3bZfGIoeyJR3nQy78
crguYFLRF2Mr/qpEkbtQO3MKwQdbAaolx6ViED9nwOkhlUaSTU/rz6IY/gnaKEht25V94hltIddG
2gbd5SwFAxzN+joH0L/hkIK9TXziHKaOPR4sOTIAvPolKMhe2aFm4l/psFsnEWiTbd7oBrb7WAHa
li/pTrk7BO7UOFgS79GW2r4MGggNEnbAHthN+fM1MOZgrblV8NThm9/jXteFVYYzT6iVJpHoPbs1
2R3ZLHvdLEeftfmX1vcgN8HL+HRm27IZTwkR5JRxyIjHep1/sCjhNklVh+ffXHk+MG45ckv9eBz1
+wpNik8hoYoam8V68gZzKf6s6XA5J7pHlZTl6y1+cg4H+FvBvm33cxlUin8usps+OrsxrHNXm05k
DwfVLYeVGjNz891YQcdedrWZYJqDEKBv62T/XLsVYWkwJDn2fIgF454MXcoJlRhAGPg86b4dbYnA
HR3cxGZND6P5xIdSgD08By69DXuaxDhhY3fAXDJA78FP0NcfNyhwG7bz33kXeiIU/eye+75XWzyL
+ZSgUtiLariGSDhua4xsbgVSrx+z158b8/80acsSNDaVO/GQZvV35i7yBoimRpw3gM+z6GPH5o0C
otqzmmjic+Bjq2bqyWvK9nLOK+rFdEgkSjVLmIdJe1b6TplM8GSYMs1IGrbNGL//4BZwNbck7LWu
2u8R8EEWk4YopwFk6TGhI/h89VyM64kCu415nnK2SuZtrI6+2zZtbHkbHwOHMw+v8jsOBPf1MBeh
rpKks7akFP/hKbJ3p+0hBjDHSmCkfCFc8n97LEkPzuVNixaeQ2cPKg6n+Y+fnHVPmd2Fp27iuZpt
A08yO0Pn+lPVCRZqA7+lXt5yNGUxfd+7giTnOHFrSqgRPLyosQ0MTb6c5fPifUjLh2Hp+9psJLJZ
gZFmT0FrISL71oaeo7c3jQFQSyVxRFP0ObViCsAMzOyEMqHksM7wXdaQE5DTEnxAS8fYEQ9DBDSb
8jHKU1/TNiaAK2tRas0Mhi+UR1FZa6uSv+A0mehMT8AJbtkFQrZ0mKi46xqBSov4UrktUnK8yBqL
iW8SkMRua9M/A3oPpz3hEB1AkiMsGMsUTUKO8uqVnWvNCSXiP00Ur2kBYb/Kd+2o1eN1lp4Wt5Fs
7HqiY+0tGfoYbxP8NZ13rNV7/aXbpnZHZi8GVyoawV3sgRAe45+20zF+NUC5wSnsCVRGdTrlXATA
xEHjdT/O7q3N4LXtYFo5B6XNrgSIrRkQxTJGLr1lJcCr23oLrJyPzhKcj3jx4Ft+OaZVmcAAM6ej
P6VimYjSHHgwu0J/fVtow0tVBHeVh6jUbumOExVnQRdkOg0jI3w5PaKquG4bme0BNzB52VlwhR/3
TIFKgoZwxubAUYdv/xe7/mQ53px/ITB8QdZpMrdY9/aXZtbd5G4Rej+oD1+IBoCc10E8oXXdywRd
jho8BA+D9++bbo6Z9e56rdBJsgMNb9G1fzT6VEFM+ngEnvlCoZq04Wpi8sbchLr7xBAmCH2sDXFc
R/gmeQ8eA63HrIhxWfGkFDGdSAfUUqsif9q9P2mWtcsL9I4gEZDyQiFhlTNHDqw+r4be6A/YSGcC
z8eeI0qdrvh6ffaAPrjRSwQR2PDkgsJeQFLGS6etQgdXPt2LIl+XS26+dKwWQejhorZrhS+ZLgYC
YSzJxROkEG4QeviGU1KrNgMqB+wLRnvu2PbrAcU2LKrdmt9EXSueDxaSuDhzgG2N6BjR5vknZpMA
AbSfku63LrAFQLBpElmU4SHlI7pNIDo20MBG/M6Gq+xluJITtw4Gk50964FSl3bERHlU+8W+UM2n
/Y9TbSNKjkHK+cUXSij4CqgE4jmoZ4q1qJyDsXZd8FzUKdEH2DI+NWTuJfmpfkUePdkIauQ/kr/o
ZrA80bt+Y3SYTVUdPmFcOvW7Mz5dYW42fbsxenba2c1W0AbLjHXBvvaKXY3lqVqQdVVLuy9k2a98
/CzGe/l+fmMT4OAkAn8m0rXSRf8NVopXNoTcqMBJfKrZ2bPOl5g5t8Tcg+9/wTe2Rfo96C88LreM
849qUjb37WvZTYh6KKZideOxVu7dViZBfm5uOrG3JxM9lN1YBSpKVyJ8/gVy4HtDWEs+fValCaV2
+J9UNSZg419bS2eyapbNVtDoGegARdoIAbgCZOCiNV2MjF8VDk6p6x6p+gqj+pszfjCfu4SXWEan
ebU7TESjtAInlj+CuuqdNb5GLUU8+aGfR8heC2uGK8FdP2PjTCaOK3YsHrnclZL8nz6zxdJ1K2PY
lvkv84UaGr6qiee4YaS0eY0tUYXPfCSchIG14M4f8wi6GUhNZ+f10MjNbyX/nVBlk89pbn2KTYaT
wx1D37fS57V4e3yW9YbsfHZVwO7yUX50zSEeqDdCihfB9izBgOh8xgQwv3779M40YBFjxv27agtb
m5awhhjmkGB41oiUhOELfRQQrFn2vQgmRB/3B9GZoEXyYXUnXCvkJX/r8i2FDfpyPEKMXSLmiTj7
kSs9jcXz5PAVicLw+otFQTxzy1kyZaQbRnFFnYE+0hVWj4KFNAr++ocnQJvAhcVMtKDp12105kF1
yI9hikDzHivSoG3SSjCV8LzZFy7rtsamdFUr+DI4l1nzOhLwfY6GhFKpxiTwYgPCyM1OOAvW8GvG
SJHNxnXTDnMvBJE+m2NCf+IOD/3mm2y5LXFdRvzvSw45tJYCGY2Ff4pwV4ULr7GZORJR6dQpzTCG
CV17WrSxbRpCYSi68gG4UjQPngErmP+L6FRfTcumO1Nm2EJXJx7IyeiKZ0FgkwXy8T1d4pAFQOep
cQEQ5mvEQbxcYRPtQC72iOoGW7t013VlxnP+PwLFov7Rfnn6yltVtWspxgtrji3iXSz6XSWUN7gt
0pCkDAX61i21UgkTKCHYEN9YgsigG6l4AXnc8WzJ7hrauKsGluZuTsQW6NR8mKLf4dc5QLqHi1UZ
0B1D2Puw1S5dn4/bHIpyLzJg9rZp+MphO+itWQRkZMINvnCLTv8OLxfm3CPmhcf5RD08IiO7n91M
MdWZJnsiFjtHfnXUtQBig1fRu9FpCw8XaE/e5WcvqpwtggbfXClRgnQ5UJTUuQrBhwBfmD31S798
ARcS+nXX2jJFy78YFEM1BGdelJBesdQ1l0/s//6Q7p4U5mUalrvQIf3KnYu0/LlYl+KRiBSzatgz
b57HGCXzMD6BjTVojf1EqrMb6tnq2qmv6R1ufO3klxludXL8L045fXvLjYmAE+h4jXfP5GKGI5Cg
iwSf52/K5TwY3wYEccey4YvfdjQ6u8RrGOfbeMCIJe9p6VEn5v8ee2hy2NBHo4SJbFC034g+Bdix
Ec65Zf4gBYNGRG2IPa+YP8XNoTdkAAJjeLG6Bve2y1hEXQctFROaIleCw5tXlhC/MjGVwg784CUU
ASNuMqJj4SWUVW7Gjhrsx4SomS0npn4HDxUkoBWfA4DB27+4JdiDdTNOHQMkFlHth1+U8pYlOXtI
qVcf2IeY/OdSKSyKzc3WluPt204ls92Tjwztzsb5ucxx5CrV76yOjeTL0KBfuGxLK2WNpBpBWWlW
ZHKjM+nC1iUPgaAduxTfLcqnnsTqYvO4nQWk2kBq0ikHBuoavB2tg/YgVPC4Vi1gU+UOirUaSHns
HXLLO8GKCVOUzLuXahfpr9RufTItRc+eTjetAoxUQoK35xBGpBel9+Of2iLP6qh+s1tl8zCfzOtt
aN14fGKpg5Fkt3cERBUMSnXnHtKNv94gJDFiPweuG1Li/p1Lbv3yyu8IlHmJlUmcv4JP2ENajifA
kKhdG5bSMjQbGG0Y3EypPZfKLSvXZKa7PXI+2oCHJM2PQi175EbyqCQ2/WxMjTA5Pxbge8+4/dCw
wbCp8RdpGPj82EoZfMDiWtIOF+M9sQroGvUL26+yyx7lDS8zUE2UgXvrxaOvrWE4UQNMKl9wzlOg
3PnlraHqZL3Oxyh48mAoP8dgsm6fB6z+221BNSjU0leZJEF7m4B8NzZqm4lamLbyCfGyQMxpqRpW
hTrnr+OTxcp3owqXyEzJeHxfw+EBiOTxBc64sEL4mBf/4KYmDWDcAX8MzqEFzfUB1XJ7s0z8n8ZC
E4tW1FZ4Wn7D0H77fu8TrWmHjCq4+18E3EeBk5KtnbAmkF0JKsf1A3ODs9kbd4zqlzVbV/+KFvKy
dMFmjxjkUSEk53wS7Ns85ujlRiiPr6aJfoxK4t4Wv2zp+2m0WNW3ckMq96OhcfgBZBI/phYh31s7
BK82gvAMK2LdjoohZdw2w9Ak+iHb6ZorAvdc77Dw6w8bqdlJZpfN/I+OwX3CtOvNsRGlzXnMTKNO
U8pThOOG9P96L/88IrWOXmZtl6uYd1gQ2RkQdzNiB6RxDnDMpgZC8aV1PkXf/XXWMoY0MZyAv9Zs
sElEba3414xHMGku4KhjdE/Rti96Fsryl5FHX//vQPuIZZIogIBod1tDM6i7ngxfmKjEBbW/DOJj
8GDgocDkxMxMJPB2xQbMuvty74ebE8/npPs8LWdENfyQlywDVm4DuRHkCUVOuLN0rymZuGR9puno
qCR7Hb8alURkFQd6Z/QK6CYqUau2pRESZtC4KEwLYw4lP5roKJEhhiFwlYBNfCqsak/hr6kLfeWv
le6ZmSX699wz0Oo7Ie692rDw5I/LPnavC1qp4/5RZM67hG3+gG5DWAFP7IcBiLwPFunGbc5MY2ca
QfKjgHBv3oYIAEfLQaguffgit4xKZDBG1C6MuGVT8HNAVhcvt7vnlGPh4+WmAPfv3femDN/Vm4fq
/O2k+vvc9+O1oejErE2lP/xBjT+PGffkGSTjR2Q4JKrEFp4EiujJfOkZu4I0dwwTEm884UkfcgKS
UozFaPue5f3+62EPkxCqHO0w/y5a+yb+Sgl7xMxafqv2VpPm8NJelxDZ4sxGO+2ON9+phc08Oli2
HHqyfEx+uNNu+Uz5Xbo4FQ5iXasNy3QuXfykFyPknJ3D721xkSg4xnggIsWcijAc1hmPpCR6qtL1
oX43HXv6A+mPxxb4urJUoDwIPr1f6gncRaCH7Isd1tHjOozFSuEi5L1/T5NdshuIEP1maR8rkg03
rnCvk8j3MGAywRAj0SjHIQJgKqzjPWH1G9NV2/GPKSgrYfTcMzxxww2Ndx+bZebF/QzRcvv2lUPY
Xws8lpU1eA/o0/1/FFJTR+FxyJCnK40Cr0i5VOllTh0cj51DzOCdOUVuLL+AOg1fcM4Je+Fmbuep
wNEuUgMvXnVLSLeb9FsopumtL0qC22Ct5iCEH6Cu3+dY+CacqcKIFhK7tng+uSzbLp7emFIiewQD
dfawyEUBpYfVruYeWVqXqnwTnKDI0McHFAuZNHXkzuoAHYpemYioBuzxciWJThDZ36beuJVELWbg
YRskSyPLYkqbrnBWns7lMZM3KvpgEiAEzyliLX3Z5vNamOMPvQt7CFr8rM/0xZL1mv1DA68Xn9pB
OTjNyaWTFOMQgdrhS1+dpIAHxbkPsI0xd81+uGv2oMqKyZ97OXoFgp7oB2a/GzQ35Z2TXiw+nlMv
7Cl3ADwtvqO0HIFSFdRnN8P1fm+dmWmiZIh5I91wUIkDs3mU/EEK1nCwYFy05pB25JjqyG9tyrKX
SnXc9ETUbac53eiifc9TMQ+OYYK8+kf++hhj8orJGHbU4W1Dew1qfV1H0+NHGfefRZofuPMOi5mC
rq9lvodkkl4N+oMGTaV2qlBgI5HCZof/cB+fFlGT9fM72k1Z9snq02ugIMrfQugBfWlWt1V402J3
3/CAcmKclliypvQZLbLdnFjAwuTb3QFWAgn14bppe4r0rbekcNPI8XeUJSmt38TbyOlPNdpiEWkG
Ho5TWWKI0b27gaJ6PmJc64CmuPssKuxb+MN3LS9gK2Y8qMjZzteRvy4CBOWEQZfc4IDHAQIv/lj0
ru1SGBfUwQ7LYOjMgQJn9KaMvts0ZEqKaC3LFKupP6NjkPEarSTooI+UmGWcXI3lGrJZR/nv+Xqa
TA52enRss7dZFdEMduuN9Y3OmPa9JGygeN8eZ4M25cU3N0HBIkjEEYrY6pswyIeqHrIKt/X8AqB1
IgrwmePk5o3thJ0nneWDlMz5DCMLj6QxKnIsfOggLK+5/ClYSC3eeNXFmfLPskcTBNJPNh8wrMen
ejh2+P3mDffapiaX14HRgPaAveL/2XCRVPQeOSFrVropvyFt/GK9zyMFHa2+mKj01zq618wcQCAh
5n1RdPPFKdyhOmjgQJnFhbRmsgj0Q8i4bG8Qcfkuk3QzxLDnECMldKgqwApCXOhkcf7odFaNEtpj
bYcU3JBZGx4oGmeoXWkYQZnhy6lECMPqzqX5GTzd2Q5VuNv9uxLZXDSGVUuemOw+xSmjNexRW8EP
04khDXdQVdlrkvtHYhBWfEyG2UimXyYlXVR/ayF4bt27rr4Ce4yovcUWvqZtQQSxcwOdsL1DxGfC
tijWakgy6ib170ikMf7KvRgSQildM5ah8EJXdccWQxN+tqdq92u8p0UQ5OnBw1uif94HIM7vtWUy
2eg/pWGMaKVIba35u+xUEjBD87hJFctHZtFmIg+q+cCbY5XL+rb33rVJHAuP/r3J/7nBK+xdbpQ9
jgcxoIkNLIw9haacqxLTYMdKJl+vdeZxWyaVZdbYAo52ssduZfL4rGxXCgZkja7xukEcVza4IM0+
ygH1+D8xcCVJHFQFj5HS3BtHM5bpvdAjdfJa+IzvBoug8nC8Bk1kzG3xPYxSpS07cG3XyaTQUX0X
BLvezNWbF8d85N8xYBoQvqJHzh1y5xZ0hjSMz9b4ldwdQ+7Pmdji70hVxwFtwJPb67OW82Drrzle
/V3UP+9GlPUdxAV2d2HJ6UVUjY2qvjki9HoZKCu1mvBV9spoD+BQv+iqrlahL/71tQ8N0ldx+zrt
Dw1fvzulqo7gh3NdWjONo93rF87ihMgn0uI961IlpVZtk3+yIUbCfWA5y3VZ9z/x1GrgwLEgCuez
GYoDIWRXXADdxr91c7Rzf02AQLJdgNqU6EkiPSKyX0yD3dcsvH5XpOXEcPWuZFfn0PnVNMuPLH+P
KNCUyfX2lB8laQHk0nHftq+fAIh6dNpit5ta+wiZJ6ECCFC3gPnUorI9Yr0lgUIWX4NJ9QJDfVjg
s/Q49zU0974zS2g19D/7SKmStm/gAOyrhnWt7DuMzcdKjvb2hCGv5BJCfkqdr807dSWVoOz8cH1i
IYJ4r+eLHtpJjmYCM3I4oriy4y5+n3JjXU49PsQjlkkVYcWaoOQ2wYXOKZuvGxQD4UTfyzlixFW+
96XmFGr1WVV73EoCusVzhZElHAO/Tfa/MR1vrP5jr08JL/Li0bOoCT65rNC+AODrkZ24NfDbm+P2
wvWPSpk8gcQkYaYrXTzQ8yGrBo5JVlCLOljWR1Azq3jb5QyKhm4MdDa47Z4CMkL11vDrsDi52thV
p12sqhtfgtDmpNZaR1LtVbjnW+cwfj/RJIihisxohPFXVuq7mhVnr0eCUYvPCyl8GkrDcIwLNYvJ
p49HbumSKYGSa7lonFZmttRI2wusV/rTKLa/xWTCZJQY7KM4nhjAsjb72fXG7TpxYUZVolJcN3gy
3srckVu1rRNd+Y31i2krAKtD1vssBIvkF5Yfptujs5uLbT+eBMaCRe4vie5jfcsT1rHzMtfCF405
gFM/PHbFT5reKW5AWQ6LD180Veg4WW4oWbeT7MZf3siIIdFvXpcHUpnbzuf34tYTHIsVHNP48aQO
bHa3jSIgHI6EgGGVklnx8PfYJ10j/rhqNcBDtG55yGddY0ksQ3vRK9+AhzG1INqhgjlksboU6A6/
Jv0l6cABHeLMJlmk7fUJEoDM97yTxTfo138lfF0BJEFsl9myIVUxz6y9gEDM5FzEfwaeuzcbogTy
fr+fCsJd9G0Q2BafJDRqeb2hhPrT4C5pwju9fTRAMvxApwcpcYCIyAa39Luvz8VmtR89VDeRKxTM
QkbaTl0fwwK0JhSxiLPFlyz9lVjb+AQSXMIUP77UZ2OHZg5wwDaT5rNp5CDJ7cMSBOBxFl3D13m6
qG3WS/Ov44kwEg5wXBfcTmNMi5IbkGtlv2Gsg76N7Otcht7JsbrL49sIvXE/nwXYo1A+WCWm79nH
rP2qhQPwuTF03VfZiI119cJmCbV2V5rDTfgGo+GKp6HCr7qHMJRXGq1R7sfZm1CCHTG3YwNroOyw
rpt7OJLFuqwb0nzjBzhAyCGsqhYkhIK7+4AdzHk/+fj1HFcQktHlO38IwSN5FVhH1YfiPrIj2gdH
GQ4P7p5yQDspcV/V2G4kWLn+y5AFuLZh/TaG/L767t2eOf3e/5PonXt37fFKlf6k+sxsswDA0oC5
133Y1FXwil/601xmuPE26wc9yj35udatB1/xfV4pIhSKrY/8JMQsVBeBn9nKOtBRIwIPhk3vhzis
jviox+rXA0fpaE347Vw6OHeDdRzpdARuOyB2RzX58cgr5y8uj3doXTY7HVqov/iAWhpFTsLR/wrY
d2bloMYrw3G36xUglHhdBivB1kwJyYAyLMo5VjOWY9XhET35/xgr/Xr4vKQQRr3oS7T5zfNbnw8y
Cq5xTjclmWwh3eskMKbfmifEqR+dMujEBDTFDex5W9aPGGANWrszJCmC8UZVhQAgw0tQGu4Nib8t
3OLuyRUn4vPeFTgPDREog6AufahuBqC6YG6eJqrcMGm3Bm21pmz/lDH3smI3wfKsYAoA0/WWcvyS
V6ulK9zY8AyvHfyUmHqriT4eMiSu/NcoSbWZIN1Noa2fxUtKDRMhZgVsejPN1qdEzG6HD1li+Xxf
Hf64oils415/INR+uQzxfUWJ1VhKB9GqAlu53XqK7218kz2rj6ThmHnod2O86xJTsCYr4DO01Zll
T7Kt+yvAUvZUSL7tQjLL02aJzdgpcAHX/+0ndB1CrZWBJYeeksd0Y+qJhqHhI3ywm4tjMlGcL/3M
0gIitSEJ6nbsTgu68D4NYld/JwjJR12TLd5VJ91cOSHcKvwrgK1r/tWeuVK3efSVC/wuIBnqhySX
S1MJbvzVoCmwleuKJcqT0XVSCtAKWspGvFY7sGyv3coCvms3WFk8pIFJs7aXgw41Jp6GIkLjz+1k
9bPLcmXU6hspyzJfOL8yYRoVImaU3CLtEuPT4LZRdwaCYAEIsJUJ2IAZSw54IkdYG/bDC6MW9Fij
wVA6zj7d3rFRafaqnRptzMVvFmE9XJ5VT6J+a15UaID6eVl6Ck2AcpDG6B9PJt69ZIKDIgZhWGce
4DjkfUFZL8JQNdlpmiFCK35f0b5TAbvO211/lVOxs/WJaXByj4AprMzAtr8k30fXy2IffFm2MsUZ
uGHiJ2kcXQVpX/jA+lF5pMawHAiESzaY/62F7DDHc5++TUYg6N09L+QlY0djAkFID1/QeuuhS4z9
KWEy9WK9S3GpKUEmWmgWlFvAXxKTeCLkVTTL/GQxCevhmYeQCb81g7zbG+x9cMwWKaBJFdiZrI3e
mmEQs6jAws970AEh85BXnD7JNm/fei4Sr9N/CegTkX8bPPXGK4ib4EsquAvLHT/xDvkcWHLkUQQG
NiHzdRXXHpqgPwPSUGZx9izqC02inZgjBU99TPQnyMfQOHYXmuZM6alV2D9MWNLQ9RMbS1jqV0RL
4xkPlo6DKMjvU0sJVdnDXI21Hzcy0zx9+MiNKqBEOka5aRt1jX11+PGv91sDRybJ5+894WQ7I6HG
jRkni64FOACXd5VF2WbhYGKdC6iFAfk03kQWy0Vj/3aroUUVSRXjgT8d/3aEzaAVDFUxd170bmhS
Au/wu/GtEglrFjEg8Qbi7CROTgeuzwENVvQZOSNeqgn4D4xwkadNzKDYyOsFDMTEd3x4DyaD/vBq
+9EtRtJ5Wnvn44bkRS9mzpOYrEZNyIaI80NbPGj3xnYyJtAuIEj0sctg7QY1GdcrdVUhjL1xJnGA
8K9/BhFRwnd+Ir/B2DmP1yVP1wrvp3b6cxS+fu2/XMKzxU4fbQ6MqavS3VHOiWAgPqQlunpvPv7J
euUgzpOpMZi5YYMrgBWgzgOBAgz6dfk/stzgKHWPR/fVSrqo7REx3e3Sth2xOAW2giaFIPKsvvpW
gKpU0AEaUWHfKob6xbTl0MFtLXOcmScl+LkBxBFNw2YiiSSmXE0iaghxcuqR3JQtmMgAhxlP5ojx
piU1THHEkCbYB3rW69T+2octWoHU1ASNcgJa9ZhW6uDfSefAQ76G/kNxd8QkgLZkg0BxxQNJiUTb
HdQB2I/gXf4k/k+HiG3F/vgnbZ7dBKMK0Tj+ouq7J9GfNCMwlDfYFq5lAVRhXtwTE5BwSBt+frfW
VpABf6qKeE9eRCzSNzQ89qLwVxElYLd18k5yWnTU+MdVHVR1hE6QMAfrVS/yWi9gz1gZ2yutkE7u
eSJiJ+bAxCIeFw1Yw8pLDcx3bfVTogC19XLczQgGI25FJb7ADucHuGW6F1vKNtpfbTjPkTGN+FWk
kJgCXXZP7HQ3CTh5l9FfteatHMsFRREKo7MHHi3wfa2yHfRK3oVPgVL4NsYOOs/geCBmVT9t/1PV
RMU4V1/A7stoYDo1zIQEkz2zyIz+oPAzmTl+AML4mrWbj1ydunIrM/Qjg2OJyGmZLfKHUqf+hIXi
6QoNR8MfgYXO5k3vhV41cgsdVA+2b8lD+H0MRv/C/2Qigi/4EzeIS2020YvrL8IWdUV3mB2hNlI8
11Y+5LqA1h3642sxGuRJlcVx/zyOe2AbLcUlWGfbSXO8G9YIIWrBAk15BztLSA762bkaykVRQowj
E3x/ZpJbXNN17C07jukAl8xTITBBr900H1mOYFjkQAmok2SEhq9bAMTycTBe4bIsKYTwgOjIJfSe
XV9e8RsxiL6eZqZW6ZiyPjEvh0uuq7Kl8qjhv75SG6CqNZxuX8MYVqJUD/EzSjxzILqIotaScNgE
RG01WK631I6nw9YHYHvYeoB8GyPH7w5emAMdG5yByXWpOYrRjFHelVOWpJ2o2mpCF0q2Di8upMTe
2nV4fDFA4M5sTadgcA55saJuxeVb+jlBxsCO+6BgB8+UxQ1fK+M6zMJcoBSdDCmj89Jjcg48idtn
7WoQd9/VZN2iYknbVKrYP8pvvVfkARjpSc1lZfCwgCdMWIwpzgF0JsnDI/nD/CGYQejTXAHRZsIY
UJuWUuga4P3S8B+wo6owy74GiVIgV+JNc9+JaU86BURUL+E/zf9F96QxSN+AqyYFVppat9mAmznK
dfTw/teGMDwvMNJ1ou5DsBQcN48V5p0JJptbyTWrj6gQxXAaop9j8umj36sCficE17jCxXwC3Vpb
qq0FcYABBZnbUqC58z/3JIIDT+1GaStEBuNXd5Xcu5LCs8MQJP7rlR7K7hZyjCxRM0R7JEz0ukjJ
8v+XoX+qI4NyWw9pP7CiZIvWp6EQ67u04jpuHuMlybQGQNUJhO3hfF2lx64c1vyv7hAKRiTTOTkF
F3TywxuVtaLB5QpFBGu9YF57i+ZOO/ZDp41iDbeeaFnk77pgDUlW1Pz095rrGIbZ9gY8dBbRvcJR
HrtCfznEiuoIuCOMJOooa9FYh0IsJTI5CYqfp/bfYrs8nTR1VYGPmF/ryNlWAeipifccRfZ9GMKV
VCfnDKpJfSITorDVXg10amfy0tNuLR8ZoUlL0NwH3V9uWA4nnmORYCcK/h6UGGR7dCbISo5Q6XBu
aBkyFMwgIILUD2s8qTeRhSUC3q08P00io6W26DJ8aTwx9DtrskydvEbjH3vxsy33gfi/UriGa7em
w5rmlj1jsu/4oKVHKhOwqaQLaY2GscuvYRxJTX0jpM5qBLc4w+yCEkwXZyy66mtR5+Jr1I5Vk20r
t+8S3e90A7d+GuKDN/6yCPQTFOys0Ly20ZQyjQCBSGFfIsthEBM4Sbw5+HarBf1gpR/pcKCy/g88
tycAVC/wqRvzrljz3G9/mFpJALvsYnnlyJl9PSlri9eF8F4fug5KvJBSmP9536qwW35xkNszyM1n
MkkSe+Cn4FsVMUbQ2pORQXGg/Opz7iNfCVGbF5eOAKE7ZmkRukK4z4sEHTOJO2FCKB+HwRwrywy9
QGoQpcfHA21GdGbxNajH14WduI07IVhE6POmZYOqMU+262xy69I1ejx/bmxoCoUr6JrYmCRixcEn
reR0tID8ZkD3hKRNrjeNfFN9gf9/jcunknEWxnKhBvYwaACwKrsuafxeVynJ9zX2R3a8w4qy6hDj
zhuRWeef07KV9XbpS8ZWCv+aFEBPN7ffpPIWUDVpuKUdN3YCtpNeZF7L60FUqV7YY2L4T35Fj5Qt
gdG6D2s5nhNk7AMaOXIi0Y+xbTxp1NVgjztQR6muQvdZxVToK6xQ1bIf1KzqXDnkZXBkdYrMUOGh
WqxY1zo+BPYTRFQWPvzAzaE2UGMcL3oakivasS1cvaPIPvYVN0jX/R2684VK0Tfjkx6xRZpcmw32
5icX3T/FVzEMrdR4zVYFR2VF0KGWn6rWV00NkayAIxTNEzc+MYyyrCeHaAbo54z0c3DsheGyvH55
W13gFZZLre77Bq19SAToYs/zS4D/0Y2r+BjF2BuzhkNSZaboP6KHSneJqjE65nR/FnpOoBmH7US+
6bWOVj2CSaeSbSWzIjXdayiZ9ar/vWF8+4GNp8IaMQMUWwBxw/Hj5jrfzUjrj5h4kyFWDBeTq6zk
AJbmGpFoXWypZZlWnMAoZfhfFUWJ83CyD/hA4nRWSpgSVgFiHFfSbItQIK0xQDZkKtCz5zykucEL
gSFlR/VpmtFBb03PUTtK8jM3c9YAXERjA3aOEXjqorfT0wvajatYxu5ullhTtNzjzaXKkQcE0g4A
444tI29uDuNVXZ95lMa5Or6fTqFpkTOqk0C2CFODvINy95F/jZ3d0udhL0ouF3IXBhyw4w6j47cO
2TTX7MX3v5Jg/HLs03YpAKKf3G7M2VMkElkt7aA3pznzDtK14DWrR98itEs0ss8eY3u6m7t1w2Ol
ECKhFjPOt+imT0x1HWLuXDH/koyMDfuyFmhz4x7+ZcgoziKxrxJfcj9Ee7/PdKs1JSC/70MnbCgK
0nhUhm1JbJwB7e6VgsjKQii0/PDn6ksP/+T84Dq+kNYheLGX858E9dHqo8OUP/4dsyqIxZz4aBaG
1d5Q7Hexdud3eEhyZa9xUM1yJy1V/oN/a6P10y/+v0evFj7OoOmtu6i9XA5pcmFtD1JLZHig/evk
Sfp2B8y+zKrL+mtBRWk/TaZ2oxxDWLV2e0b3hhBO1Q3fSIQFGU9+unlidas1o8gV68Ij08YnHZsY
urDZLZQREcL2V3lLGhj0FoaFsVykyL4AdIM6xOPTi8QE1c0sXo/B99KQPHSyIakeFMowrozbdXjZ
Gc37ZMS7XbysEbT9SLfrWZAQONI/94ZelqmQZafOS8Zy7GIMI/X5AzP0GOwPvy75EOC3IZsB8lCW
+N1uOjsIA6qpmzoI3T/se4Gdq7DQ4NlcxeZ4WXSAypN3Hu3AT+8d8NCLiXC7tBQLWxjntbu71+++
ORuOfiSJF+UCciC0kyXxqb5EICWIf/IqETif79WzGrU7vtMtUo8U9U0hApbDfpbRn1uM50PkuX5n
isBag41n8rhjwV8wuUkz9V3xrJtcDJtmT02R39ZHzrpuZCxpZKCAFNFb7JgCKv7/LxHeDnKc7mRL
IZUMvFhR+uySv+7nQf+NPDl3Csryo9dbXCk7yqI66HiYqf6ywI24G7wAhDQH878VaupASlNChoVg
dMGv0fNY6lFGxmrDrFm+n5XCulmZG4GJgTXfR2Be/pDXG2D0A7tX6x5I7FDUgcd1zNI19aiQFVZ9
jML1Wkq0LacLmIoLfkRxUfcdXNS7dABccGp49Hl7Qd3QjNDy6L14gE145feKE4z470j3L1fRzqvL
hYYPfSGrB1a9JRat8XYxQ0RLF+xLsFTMsUCKbzHQr+45ad1uqb2x6aA/9EIyFWiRPLgq4G9DHHDI
SIJCyl9aACRwYuZeGgHCVZu4ANL0yi3icqsBMCTJNgilC/eTIsUDLtIGsJN+8D/QIdMnqCfbrgyY
JuXaLyob8cr7/XVaY/2SE8WgAWgFIXqrIp3+nXE4QyV2o56efjBb0jR1EDMi56sFVVGy1grS2jk5
KJrUgFGk0dszxxQgS//SljAneEJS5leyys+UarqYqnICBkpWXlC+3fGdlhEGhhv1SrzdMwSKelOa
pPP3E+gotMRgy+wx5CsWnSd1gEYCMtqwRkr+fVLp7T9Ezcp/e41/IeN4eM02E0k9WdYV7AQ0NFXF
GIXqEk6LIK9jNYriGdbEjiFT99nHIix//VMO9+shgtUXScqGp8XYqB+VkEaCCG1839j00VzZ377t
UXDtb1hiEElJuukOAbcjr4Gr7l+TWpBnda063TG5KZeFo3oJkf+cDmVpG4d4PbnR171i61uRXuDe
3cMXbCsPIext4uDWG7CopyUKBf+n5R+yWUcTO9bLIbY9JxYu3P14sKXe2UMjl+M/oaC9mUyUYpmE
e0rkJAuPDzxu+cfUX5FRD4mEmhaKW2511dEMtwcqGGb6jnmfi9Lzmjs4hEhLqBNrZ+QSfw1texrH
UghctI+HIP01qhguiETh+4y8pNBy6D9za5aeFUxnVDaT940oXApa1UReo0Vxq8TjGxyVRX2cIkya
AxlmqZOIcAd5LkbGBq1QjeJ+ypk+WNnia8dethBTgjA78hyzWLeIxZhahiFerzUbFRwf2006dqy6
5Lo6s9Qhdz7zn4OlBnAq8Ekn7aopKTjmDZ/Y2Gud84ilsP5AF0vxSmJXPpRT7ajT5xFViDGbKu61
TBVtcG+csqYppRLWKnzR2raj/7dJofbQVmi0Qll9TRKVXPnmflu/fj/FuHuEx+pOQmVNBlySG3x8
wqbBuxurSC9FmmC9w7yzzTqgYacaElGUIjJL4JF8qVjf72DzVp5b44w9cod3HskaK6qxuyhdMzxT
MrKLAJWN2IMBCGi2LZrKwULvDby77fvoq+/d1BQgQFTflWuzo8OvglYS0OLyEGOCEJ2X8yEVDmBJ
rTyAxpsfO4fNrPttwqM5hJf3Qd8Mz0h1xfWCiZewXNvW8IAHGFBIuimUF88e+7P5dV/HyMoR1KAz
iEiM8AQRn0KxQNA7u6LZcGYy7bmaTXE96iwgEkDs0OZznxR00rxf9+EoKKlEhsJg2B28uItMb1BM
79nk2Tt9FyRzd5K2FtdXZrhsOIUPHUG1wrN5OCkVkc0mSoWv83a2qPZD741euAvUk+DLchzcjJ6o
/490ahWM24wWMmtv1zC8K8/19xw7aI+RrmWsHyU4nOt6MHpdYjGuYg5L28lr8PAgjCZUD/ZwAUaf
SpJoEE3/hCxpCiDaYyM7d3WQUCxCap3KQAM2mXkhJSz3Y9c5kjCpqgleJAz01l0MybvP4/WVX+Hs
hhFkFIedMZrnp51+/lLaAc3Ln1xSEdcW8I1yywPKKUDQgTRtHoptA7vnxv0gkSypA+IVJMmCtcuN
n6sHlNRektGANjsHi+ctLMFX/la2NC17KY1sZOpE6iPXL7958jej+hPCDr8TQwThy+QuSHFGeXvB
XrtvFZf3EBc7LtxmlQHN6kpSpZQ/oIdLSwd8Oyt46IrKdn8+kSLm0RagIPD9wzNNE1H8zmCDaBxS
TbhGytVJhO3tuPuYdNSRsdzuAY2DPCT9K/hhISZbwh9barDMWNnZygAARrm6wkLSX4X/iF+hiI3I
sU9P5nqRAYJ5idC/G/VS+nT7O5Rs6lW/FqQeE57l4DF4AgtvcolKdYTe9utVY/yzaTKX2jKFELEe
2ZZ0bZ1C0nsULBIOoQDt0SJcxIo6j+iDVV5o0a5jh9lwinxTI9p5rT/7MiM0a5LAg6eyQSI1Yjk+
dVHS0vGu4SEOi+oqh0jE37VHF2s/oQdHZN8KL8I5UcTo8gPQju5Zd6MHNNYOZ/Pkp3mA3DDw11bq
D/jemtrFNoZJFyk/b2F5jA6+R+tZZYDjDEv2f03W3t+vmoZBUyn4rd55vYRH4jBj68osrb1kimnW
8yPCX7e7oErPQDWDBGVZGa0hR8ogyj6KwZgtGZrREjE3wrtcYW2//9iwQHxNjyG+5gPqzlS0DXWD
1hB6LLjyBXlgWvDe7rQCa+Xo5U7kp9wL10Sjf3G7H9kkpKD7CdB+ugHl27hL16+5bb24OG5gEpev
AiRaypl8+Xjd0U7X0g58sVkXaex2O1PbuS1KuIbZbJcRPNgp4JENksrhelKnRCk+3pCNPzwlAyZ1
D6dqoDnEGdI+JmBI2WHF2MmscpIqNvTmYPCSUx4khallr6tJydoiZkDDPCAmgp6SNn3AiQZybpZ2
RX1GJyKiUsWx8lfEQQf/GYk+SXpXzOfefzPObVJQ9+25smDoikIJn2tOkcQ3dSdRKuEsJpTscGFe
Lm7S9ArcruTntkAOXMGVCpS/qp1jIE6k7rRV4YHCgdo68UP8ncDwGWWC/+HjNlFpy0SClCgVOhvA
GTMoviNJk+hZS2hHmm3oiDutGA5WIiL0v4Flxy+OUYQ0iBO/UuiUhlrpu7n9/bk9t6J7AaB/hWn2
nC38jZ/Pe+IPgvcN0H/wkKx7MACZ8OKO2dSomcUVQxFxznteEcC+qbbMftEnBd2iAs0SBjPzhtxw
xQ9gDfQ7QZLwVUd63dySgA8+SgSHlclq5lJDfMCa5IGlZT8XEkmj4W9b81q2CRmCs9xzruop1Kwp
RF/4F0XxsMSZQuTr3Y5CGlFTB+fevj3Wsew9mBIoG++YjAGJs/yMSvXnLvM1PrfBE2pKEtnVvss/
AFaGXlLpPK9d5NisO3C82RtlVshqhw+cBZqcnAD3mlc10mZ3470Tffyx8oJ2ODRYO2Lwn3I+Wou2
mw41CKtuS1JreLfrV2ZyYoyWmWEonK4XihA2PsK9dSxH2/ebNQhEhtZy8BFMrAL4ajzVZPlrxyV3
uQio9HfK90kDxA/fmApwZH4MplMtRzGEwbfzyaer+KclNouRXfWmgdvNPIWlSvM0U/bV03gb0Qf2
347l9ymTMCgyz8mpDh+LvmBZa2UbK8agvJF5EML5CLONyXAgdLYJsMbWTQjLuHeQ7eNZE1KrUL7F
DbDaFcL8Fcfn935S1iwoa+qP0Y11RVtRhKljQ3XiX+XQZrxB9s1+5xFwIQSCtp1G2Mfu33tUk82D
HmMja57ZSaij/7wQN/Zye7OAKOZM8S/7KUrE+fbZfFtGmvlXQldJtz2kVJmo6IYYYLtUKaiqKYKS
nVAVSx6hHEVLZA/s2YibbKSSbxlSGW7qTlfeC67PL7kMKO1yQyMCRT7V91rFNC4Cney8xEchA8Zy
Ag0jWBvr1AgqWEEFaEaom5m2EnMK8d3WnKRUXAshnW6Ra7UjZb34b3Vg477wuVvRSCYRU7Mb4O+D
Zzjv49ZElG5vMcZs7C54iVU3/Y3wGLfwDXY9t2snoqQFXctiRaftquplWa7hwOUFFinEc5evPTw4
BWdKw9URYyzoF6Xe+sVLGx7P6zbmWpPo3h8KJzsdG5hlHUN1PdDe2pJMabnRWoBl3RLYKwjMgxAU
oX+qRYhR7Y3xV3JqaK3qIR2e4e6xqUc2PCPF7MJWupKss224vGmJOMObJZsCfOo5hsPw23LRzoqI
LQ9Oe9O+vBXG+/KEARtlETHnG94alWUDkZ/pOdeFkXJbMKVvP+iGLQijSgvevwK6JXm6N5+ws8kI
fXR76CfZz1vJ5tD9CivoN8miBQzfGMLpJU46D/7XrWLDU+HjX9CbGeeLlQR6po9KkL8egOqyM2fn
bQExMMKYdsbH43WS3g07q7cdgSUYFETgh1JP/4GPxBueBJZ+5Q2Q5qycHQvhIflKm/4kk/b1WGgi
yIsfzH9UhXyC1GHABFmC2ukXMx/lVvO9+t3e0mItvfxkORaZqokPl8EPMIEMmmdaG7alGVrsOX4r
ZhP0/L2jF7TeQURe/ghB8YmHY4i+Y/PVDue8/gzgh4/pU8Vrk++EqTdCbmR63eDbT0HCD7l5/nSm
1QfgfN7DkbP4fN1HOT2ctHu3SNXZgz0aHAfc4hale2IJi67V7zxJ8PuXJCCurt0WsZLZGf/gvvIh
92p/xvUW8twly1K87eQ+uQyjrduVFU95euqYN7sI0ZI8tlGKlQOHSCwlLPRsvAvHx4lyNpePmzTU
nwc8BLh+iPvNdNDe3IRXMkhyyOU6wJ8bL28ET6kjK+7cY8Ll2yArFtJercFuIndyBCE0cCHpGtpC
bMwHN9xXbCuPwj8KLrRIrAjiXvAEejyUYpFXP/wQhG95BArAamhNPRPM3RryVAKdT5ojOGNha1xQ
/e+/09Ev8QEr/5ecw9uCZWeHihh61EXwso+GsaaXGAnvcmY5uhInlgYqAsbvN9aeaLOdNzFUpFsC
Ua40LjoSQVR2iXHSxwWePy60l0DuMH346ThsQFLAD2gHB1AV5uSsVlBKHWS/qXvr68eGRMl9f3id
CSCZlZfy8UTtXHv1xIEuekM+I8dT9VBBwcWYTlmLhswU2RKzy7xMDaoDL9nYpTRUp41KW5DZWrKe
+5hLlJDXscvS3tVf+b+5o6jfR25jqLvU6FLRpzQeiryfXC9B5DQK3aB8skPVC0PQaFHckJLVRa5P
l9cMmBVnqi/++SqmVr5WYi0xd9sdcPmjvdDAwtvIIuBtdDK1TRixgJWWIeVI41u9fZaK+/2G8pEx
K8KilpUiEm7CTc6JMvUCZ6RJi026yzP9ij75vzNdOTdeTdAmCU9n8d4/h2LMNR/Ac0L04cMKTtNx
YNXQbxnJ4NcO0YjvixlYi6S7wBKK+ufDzMlaLxfo79x58pu3MXg+fx3KcgIPc6FrXiU4Y177FpBE
Nl8jWqbaIrvefPHVn8Z79G9GbjXiIZKryOG7emIncDv38n7sxWCo1fe/1AwVSH/cpJOuRU4ns2lD
1+l0aJCPfnrpn9r4qNHb7I4KA+ysbpk39gpIFx+b3vwqjcI0t9lokdJm4HHDLGjyHgPGgrt/YhgV
OOYSkwwmwDx78EUH/4MBqRFyOHJcci73rMVPJg+pEAvpas66HSMguB01gwSvUD7BFHix7IwF/RU7
TF/ARFnAh0fL7VRwUBUSENB7y1BoglEMk2wpPR9yvkPg3lF2VnYEGWMOuS/GRXbpZRvDuEpEjRpm
VKp+RGfW0WbBJcQypdMnI+fY5v2hMAURsAVIVshHu/QlKLlkZGx2EWMzklgBmpVxmch1IleBSXij
TCWRwsT+6cETitUsPKEcoB/uBJEMCujkvDM8lxK0kDHJpoKkIjKvntF1rSvVN64nSrfXzHabrD5Z
7qsDx1PQGySdPrjOFLf9tVkAX9liXieNgv6qBmRmKi5SFHr3s78ec+977lbX1XL9owiHoCar+V+n
a8G02Pfw0kNDACocTrOGd+DzW2aBYGJwBIuq7/rLMW9dbcMR4DLQrhQCKKowpbREjmFFrZMApvLT
Q4aqEv/Fqy4TEq5MForKx6sdOH0uh5+LlH99pKhMO3BTTzgNfIeASHdKdKj2oIuQoA7YspIdsvC9
PzOUNKd9+i+SCnfhJjpNdGU3vhVrP2DWSDhzr4ZX202zXvkWS9SrnjMhxnNMCCyiW5SqvUJr0Beg
FAtcfRlPW6nFRR+EkavJax0yU8VaOEwx4xMmn3O14Vii9/Q8fEQSYEwCt1GlZFd4kQQCKh8fUbrI
ZFMxL49hHlD3SZVrHvpfQbCyWin3PpIOH+RCv7eCxDyKGH9pbt2drPDhTpqh+3rJclufhiyrk2rC
SEAFE0+9GAjDyEExlv3mrzzACULwSikpxGhi8YUW4yz4E8xv2Nkv+r5JaAsSFeLzDGib6fNqi7V9
hTGOJa2AdvTNUJNCZtpMEgrN+uSPhDVmLdf4ip5ye1o4lyMiUafWJKWdLXkNecWPjmTOwlEZX2KM
BsJRGjS9pJOQvGz/9A22TY6TrMJvs6seMhHZOfsSwsYaWhJB2OWjwf6wbOaXc1KsiMIQN7hy41KR
j43NOMuF5Q+rs/V5KYZnAFJ3coQ4b4mH2D5C6ld3o4pgILbD++ivDhKcmFiaN0vMPcqXTzNf7E88
1DbI8DYBzgz3qlTy8aPoC+jLtcaG9l12w8kE9HZgWiT5A1FlGlX//YnMO5vGS0//0xK/ttOVSnbl
bYpicHM+R6ObKuF92HLQWW34iFtT7eIjaVHW3sVMMSs272uXRC5b60jAYIgblAP6Sib25kX9Gm9h
MuZFmc+qKHOlTrOBH8SPCFI9hC6vN2eW7a6fN4fUuqROgBbGipx3TlQ8FLXEhfFggG39rWpvNGo3
GmqcNmWKWLr0za0guzssDB8hh9lY2QhiVwMG13Z5rkPc7ipy/kZ16GEjPMfpp3BUmVFnkhfgvF/Y
2f7E7yzl8WmnIfl9czFOU9UJ2YAOF6ThdmURCezHnpbc+7hwXa9ARxJ26uFgt+k0fqqAVCNp9HAV
2iqzC+i+IpSXalEXQguDnSOaGmRhYbhw5OUYZgvR9Hqa9aL4fnZ4qpprfeIZ2/VZ+sqzdwJnLjDV
U4sQjCrLmVLG0BcH1eP+IH/UKEfFOs5wtvEe7zGPK7Op7qWhlYNxSHkYv8uyc+RgaW7E3+b9O4aq
DoEdedWtr3laNTpwQk2wQPtllbdCjwDtDiBZvSNdCyd3faOvJkDS/E+uSIFhf4hH1Pm9y80V8syP
meRKMHhcS5RDKmW39OBxHfBqiXDFVKcMMHo+gEhAp/DE/mnphQNEZ1ApYwQQhChX2t0neXUtRqk3
cdkQxRLX4Iu4QTaCL5QZrNzpEVJd+6mu7KpGUoxbKs2SGF9OzM1gCE1yVzfcHMaHMDwTfOAUCUkv
8xEsrMafxyjWbGzL4h31E80YFR9KnWj4436lJFt2q0psLsWvvdeXG9hVycRy452IgSyngb2bkSre
xzCpfFj/zl6+tgv9aIKnYVav9xWZM83omuC6Eog1fRYaqGGAf5bCMfcWijnHMOqTmgrIVvhY96zQ
bIkap0sbtIG0UC48wfy5k31w2NLNTooWAJBdknzfk7xpCIUghREfi/riVdgun1OcNkb/qtA1nX3I
m7MyRa7xxxHeK7BirWHKF2f7EnSYq4l35mdEh5QVZmgr8TeXskRnwd9DtzY1nIlQWQNV+7hXyEai
WQSY1S7iIaMkrZjZwTuTw8rdsNftVlsPQXK+iOk2BOQqkApmWpyQF4Sl7+x1pHfmhgulgBSo0Ivl
qVjCAORWpuvMiSkUYGG6Huvyf3ZDwjvZVBzABY4cROEh/C556ff9NOXVxxvKAtO9fWmMlzMUb6Iv
QD3HTMZUMLMeSUtDKmMxdiCe/wg2oycX2G+w2vmq1dQ4oX4IqCqo35nS02LTsCEJw2EeSv61ySBM
vCspWZkfXYyxkhYoVmjjHuBVV8H66JCtbMY87mfZhYOPbCuCVtPR2yMGryWxIppxYI3uTdD47Sgt
prtVylHO+jW6HXhZ/HGpIyeyGVNS2o/R3xVwyT+I58N728FknNheXszbyhhtgQbM0C26R3q0I68X
X0QJXfyzAaqkZJ+/2Lx5kQzET8dHzd7gHopE3nu3IF2YOWiRaMbEZa9w7Ergm0BMElLz9N8HvH+j
1wZWXvbvFBh2meOmoE0kN0uoStIKwspMrb+hyAa5aTCvyvmo4zk/OFz5L6Huq0yyXkIiU9RtKz0g
kEzuQas+eEK2s5U8PL+Gcs2ouU2uovIW9AszBwMf2sI1+tD2nbAFxkP8VHt8n1R9cybnxQ+6Z5XX
dJuM+PaYLe+PL3v/ATUBxGDf8lx2KBgdK5TwxFsOhxQLNOmz1pje6F/OjkwjuvJlHvqPkZNHYZX5
5zrj9l73WsROxPCWisSPjXu7kzz/qqbaKYMogKq8YnLd9Ojp000l07N2uqUgxkzdXFL6h2kkkECd
yepqa9JtO/kin2ZypxP36J9ng9OiTyE7mAm6G0fn6ZK0R2Pg6cEeF27xNdbmdA2SPqc59F84UFtd
qe2/tW8AXYw8RmFllWQ59dk1KxPkvGNzKLEsMK0aHsg/s3zp9/EYQfZ7k48mPEPkKhlXSZB4vYyX
Kmn26dY/SERArvmy4/Iu7A7sTgxar266gmSx22+BH1nkvHR2LCnRF/88xJClcrm1kn3tpn6t3S6j
Z3vmJF8eeAt95RcggWKfguQc2wC1xzCLYl1/Vb3VUkgZ4ACv0rJErbRfS/5gs8bt+lpdG4qXTvaX
csChrGp14tyPdMDGBGpHag2856n+jH8VjgOSWvl1KXHHLXEV3aKQtdOoxn5HSOUCQ/ojgKsy/ajT
/tIA9LDY8f7MZmCuN0rn00x47EjnAmyxq4jk2B9uujV3GhYdD5So+Nu/3sWTTvShSwME2Lh6o9ii
QmYMBvcAqphTwMEjY5c/1h2TrFVVhWDVVFD3XIgDFV1Cxtx9q0b6KdN3PgMxwp6MIh34g/Sxvmd7
WN9+GGVsPWSyp8aysbzOaU5WEckzGCp9M6sT5JDhS9L/UpfnypcMKIxP5OcxUcPH7IWfg39KwxSK
0SMrHvqP5yipGSLVzE9nVrUUe0cVS9iTeVxHPWp+99BR+Jdgq8OY2AkxCyqZIWeelZlvTws1xJ8K
hCGHJhjjgvI2B4S4f6f9LQFD7CtsW4ru+sPFTBTo9P+JcuSqJcewvGZ0Lx4G+BTxRzWtoY0E4nF7
Znex4mAkysvQNFh0ysv/j09OcYQqbzgHHMLkUsomM2kU+lBtt3u7CG2GI6qLbHdE/QdV2OJIdEiJ
PotgogPE2oDbu42Xfbd3iugiEAU5FNk8Ze1OnYq1vOaYTxUEy6bNLxyD8tN9pAB82gaVz4kbA8vt
8qC1AKeKOAgYdLhfIa0jsFTJLwob6VkSAp6vMANbnRAJg6eu2nYnnCB5fBJq0pHlFwgp+hj/ng7Y
mXtGSDEP/F3je7P2pNz+n0mbpp5avi4Ykr7VgXFyB4mzgOx3yDOoz6g1n8h9XDN87wzBOO8hK9En
ZTn88Uk04UPszIAbY4z9fJet+pbhixaX72XQ1VG2zggX35iFIyxHmYO8xcBYsM+k9lEFhCxWLEhF
/o9N/+t6/OJ7ESpvThwESr++NRsv196aOBC1ChYs+g0atwUZx5821RkArOA7GV8pr75SyIphuPMB
JEkyTRRmq3hOg/lTsg4FRATIGIopGzpoXQgJFka+1NOv/hDbIepW4Zg/BDAL3OxFG1SXSzm+WtdV
2Jh2kH6cohHawG1md6C19oGra2xCMKb+z3FH8XOshq1ewY7UEMQ1BQ/xYS8SxYRh/PW2imowo9vk
w8VQtaRTXpUdb2MbALYFh1um2gJQaeyem/2MrkQu2tsRGnygRHJJH6LfazmI1UwYNQvBoP4BMZCI
47TIwR+Lt9NMKC8bFRIuZrVr2wdx6C05glHK0o0ZUDm8W2dbZZSAf7XqITT01ETeBRoWZANEB8g3
NHSxZEr/EuStJLw9gC5v+por5whTyi7ITANiRDIEHiQqyANr3nNqOJksq6eQkVC2n3tv1cSF23D+
CJx3+Qfu2GyWHMmz1aNJCbSHUnUuI1ccBNalU5ZqsKhLD3gR03L5IUnDQljXQwyd+zShpQtwVuLI
bxPQGhMSJZ0YOq2tW4NShRksLNNb04Dz6BBSBfIs8VmRgNwzWCx7dIXY2ZOQ0R2D0DJ8L4h2P7kU
41UA+JTVnh7pYruK/PG+ExnZVA1uCDfwojuuXQEEmCJNhHINuOor/rQtxTxWxXZo0UKp8WDOIyEB
u60zJ7yaWP4bu9Wdq60aAR8sgtHB/+5c40Nu5NMEtCQwKSE1ZaM5/anoDlt+Z6dE2HWBp2frnOAZ
J6CiwCklAnMNG6/1ikkzSDfbXywq3TCGcrG0/VHsoqGeiBIeqF1DRijPfQiaVY0WMEENlF8U5UB6
jajwwrZY9WCrii3IFajSXU6lGCVi9QzUBk8CeGSiS8UliWGKNQu8kYW7PTLLG0vXHXIxsWAN59ah
JDomOk9CSQ3LJ8rhKT/f4rXdH2YaW3p0AV6PPvd/lEyKO2xNzRWSuzCB4o0sOrTIkUbfiyWNQf6P
o4lOIk8b8P+A4jma0QXXvOIEHctpIi7FS0Mg4G2pBSrxzNElNCGkPDPHwG0YFuiusyPeKf5Emwis
yEpA3Ao3sJfNFskUE7b8GqB3BZnPD3Id7TNrTc3m4nG8BR/zJ5ruRBnsMlw8tvS9FLIWxfdtE4mj
0CkHsLs+CfcTuMLZmyWh6ZNS+BqkCgK4u/qU+LtZq+7JShNhZ2/qC4AGHpA+FPJGn8+vElCLfmjC
O+tvwoS8I2JvCQRpuTpAm7v7hZI5c63KEIIRsvCR+EV/ZRtWhfmescH9UlVaAatPRE51jIxsbp6n
g8Hftd29g7oi7QrdYVhsA+gtF+J7kufCwnkvepCA1VKTZ1HdpI51C9S/R9muaQ0nkYAueppAIC9l
Ko0B+zEbn0m06tSYe3EEZ2OLazcqbsi2lnpw0M27yAS43l3+DSY4ze+jWRYSQ6XsBiMd16w/Fv27
mMD9POf2H7i+sKkJcGwYOouF8qhbG1KQs5dXOjyv9rtafhiPHDijzPAte/ROz1LLQGgBVWwTZ2CX
+xBv7oBHYkE1I5tWx+Gk2Ghc64gQmXLkh1rCITsAbCMc5x4Heb0r3OPHXguANLbNb/ApQ7BZD2vH
3v4P0bP4GkC5uW3UxPHoVtWgNpyNLoUdWoejuMVzSFVSvRtmUsdEIagnK7mzUYTlFoOr1dUyzqpt
D2ey2IbkrtT9v4XijVUGudQwVmMvDVaHvlJcBOFzWQ4vzEEfKJI2FbmD/HsmW28JTnshg1Y4aRyt
qYjle76NERAj3G+71jbEpdWVrN3M0/ql16YV9NfIxlo2LmSC4t4a2HsiN/AnQBu7PYwsjqSMqUXu
ljdWhNDmFvmOgjnNLWPBfSqLKPMLbmxFCqZ0w4FmTlleGUwbMiuzD2tpGqSLvZ/N9dYkWPlkOAaS
EmcqfwRrQDhnE/cWWCPAszxM9m5JO4BfqSb7937BxzcBkySlh5vSq8WS+nZYMm72wjd/eXiLNNsK
xDlikmIzPJyXk72uPC2CpUkTuWAAE/AZnFDYUBZ5DUW9oD0nMpNH/UYMPIWNgshXgZmuIL4uGzjc
EwIV3txQpZqUrpKbf1WVYs12nixhuOxOsM/ApkVa0zdrgfE0hzcXU3nJH3JT+/pwJlsPn4jaMZH9
iSKBidOdnvIksg52joeEOeKr/rd1dN5GToAxBZfalpM4Ub4yNh9eUmqPZxPWDAKPqEAQkCJgwI8h
HzOtx0qcsDBiKXkaBJFhGasRpc6zjqwLXe8w/D114FKXJJkPxU1eUkX76HkxT6vTXvO6cI6sblWw
t14HNXdsThAkpLd2zb7/wvvnMqa4Y13SeBzahqOOgTHaB65CEkkqc6ZGnd7VWxPph+Z9PEJHMV62
TNwLGLwcUOuX6AmMTSBSY5Wsjx9xL8lcI7bICb7+qISBEANchR/VB6DWuBAkcdydHnYzyydC60fi
SIAPEyqXQB9Alr4aT4AA+OkIW+KXT53YwRysYpV6eBLKTYLLb0I6mMfJdhiPVSpsf6nQCjU+Q1nI
KV/NVUnURSFAX0vIJA05KgFoyK4zwzsIxHA5tsElrdMU0kUBf+6MEqsnot20eIHZbzAEha0giJmn
7orQjzAmqwcw+J1UMsT1ykhyEDLRl49v+7rOrLrOhpdZdWY3Ixmg8g5xSUGKmqFMqlF0KuXMpNI2
aQsZ6katfvo+gTUVsq3i61qA5zM6YEEpjmMp6DMq1DFaMxmoQbVjaR+zsNE7dKrsD0mzYbPKObeb
s/NgYg/pZ6mat0KxiuV06V+PDr4nzPm1I2PEC7nwOkpQUUHkZZ93B92xzf9uoUa3OuOdck+Nbjgo
EUrV1BEMFH6sW4PO69786+Z78P4nqN+H6YpLjtq6VUzuBP5Mq43EC4C7QtqejSzO+IbHoWiiuGuk
Wbko9k96/mJkLfXDPj5g/5wpdVpEeDv45neq7yoqNQn0WLKl3Pzo8FnaDMYqu0KXL/5hzzA//e3Z
Xy5ygFElasF88AH/6D5DS/pKntfbA0VSc8pjIKeVdMNgYsNLurykyxKAWB9cZLVIk2YqcXzeKxQf
MgQTbPEx6fGLN6mrLm3PWYMJNTJvEUidWwncuPfokjNTd2feMW+iJGsG+rDhwsa6dDOwnGh4U32x
WePGyiQaJA5Gl9QghxcUM1kE9wLXnJ06Pe0w7yGscemTDiPukKUs60Sv4IRLTLHw3JTfbX+eXy0p
WAY9OaRv/I/nn0TBsf7smWBpkxylqH/tVR5tbjJTpf4N6vyy3gO/n2HmYOX7i2bCyNK7E+LcuaUV
IrBhiMZU9Aw4b/j8S8c5qcjnE+1/rSU1IZgX6UXb5B1eo3NF45kK9b9uktIcYa62BOHI+nxtuj0y
9jM/EdNWeXGM4Vn4BzGufZn8pBL30gmfV396ubJDI5vxOma3v3QZ4TJAX9D2PnYjGJYPdfA+bbHY
SoL4IHYYsiAjcBTr0oW3ilobIGO1td+IVQIO2QgHo8BJaTPyQHB5QLGJ9b9FHn6pTayqitGvHsvU
dVOIlmdzNkYmslQdAvvW0RScVcWyCksvnKO8BSEF38uZoBRJyXoh5kK14wVNK+EQEvGG45/Uu0J9
eGGKqdjoojqxk7jGae/+2yYXRlW4kGGlEsdJ2mFWH35lD9CtbdQk6Fkhp+3eL/9ZacWCn4JlOTSs
6WrfL01LDseoC/00LDdxcGpYYNjsaHnQ0GiC8i69nWCbAz2iOAXmYwXPyXbpzC/jZsoK5fWDT/uq
bfo2aATLg55lMYFLpMlH3hxKiZ3vKVcmq7LmG9cuf0gc83rwt6wlUEprG9pf6GfMpA2iT8Azrxzf
ZigKR684WooEUhNyUDrAAQFv+36QC7Rm+Ue8PwVbmt7JVFzgmP2wdgdmmVxXII+nCEjY/SK/PbNG
o0kpa35exTMCTkJ9fPpi+OpfEcvaTPA+/4xlMyILG/TLH91eKaqLP/f9mq3yWt5JkFHYRFsWtM5T
BzYRNC8NT02UTVRgTv6Ipcp8+IFjOXDyBhZAu+Z9Lr9iqWInAcgECa4DxPhuqGBVDouG19Kj/882
npNeJx/Zgi4ZgLreWPKY1wNNc44GSSFxVGlYFyhRfQHR83gPsXu3QbIMMz/gzzgrYmUJbkLW4bkG
aXAMPkWKXWQmdOdKng6YNmEimnNiD/bkKonJWaR6lv353/Gjs0qMlLUgFDjZrl3zaPVBo9cFmoaM
DzhqDiC2olrpY8XfkTcuqAGPuicQNQoPgnvJ3wOuFHtaiEi1/xG8yWVyIGU+IkDPAw0HP4wok0Ue
htVAAdPzT4UvewKc1x5ywkVLoX5HXLLlq8qEbKErUaZa1tJ70adzQl4o++u6iMiPsFVOEWljaggj
9wu7eHa35ncuA22kmtiuTCOPHtb25GCb3XvCUQtvzi5G1erHomK7g3ixEeKpEb8Z/6zvDF550bdx
i9dC+WTkjDezgzcufFp4b08mcRl7j6ZjGEfq7yIeg/E/RWuyUWpUiM3i6QUQEDYrqxgkXWD2QfYv
IL2ZI064Kku9me4e1b1iyhZoiWnh5BKT4LsXdjjL13Ih6CNNvN8vch3H9Li/93PZ+QS1lXVGyFJr
BNTesxf+UaYF3shIob5/v7M/E6/1KAqGGiONDRtepIri/J99qshCE61xSprjDmHimJWwKB6q768f
tpk4romeEmKO2sg7+e97MFejzloSupIGQLESJfExQ/XkIkVZr1SD6eFkKgVAXDwBIFEAxeBcb0O4
StT/EVRzDIChpGuw09cCTHwfraQRwIjujaClLVGuZf5Tr7HFeAc08hSJcBIg5owk22qKP+9L0sx8
XojVV3rkTMf54RnIvvV/j8hUzZ7ECQ1xhql2/XhnMijaE3GzI/LpVOE4bgjh2x/4MJ8ZcRqzB8mr
+J4tSBrYa05MVI5jLUREz+3jQZMhDhrl4q+FUXgSGsdy4jYxpRgT5ed5fohrmBU4zuxSKAY0uGJY
VU5xyAEIIbgL2qoefz0Panm84xp1Pexs/aA3VhUs6QErLHOVhjjNHTyEAWWlwdeDo4nmRVCiOHpE
snQANZwd9q+VOR+9PBU7bs1Fk4YysZaKX7HHCDHVB5qG1gVH4Iw3UN/SydHwTqbpa0bhIEMhyfdj
pd0S2lzLxELtpOcNgLjNzXEbFES2Fy05Y9S0sY1tUNnq3sOAgj1tCVwqr8wCh1SaVfHmfqHxy/Vd
Vo2Fyzar4EVEUvRPk8zCgQ1EIZ5q5fwxgq1VlOzy2ZhDH6ALn8F+mIg7P7GGp+b6GsQpRHVdTyRn
nc/6QhIjLkVF9KyWjI1Kh277S9afqDy34lGTyvxuVVraYorfeehEig1rT0CIIVZ0nHJzwh8YEr7J
JW6w4Ga5iWl8KmZVGRJgjMVP1itnW1Qbjn4rbAUmSdJcL3CEqOvFVppGjRLwrnrp0jTeSiRCNPn4
11aB4gZxz18odZLsbmjR0lb1uE1XSmA62pOUHTi3Kcj86e46j/QsKwwEalw/C/mUoDLUynKWGkl5
OtkFcBiY1v4x2dJvj2tTmANLgVNR1+Xk5UR7dN0f85a6PSXPQ64yCQQUweawVHgfAcaxYweQ4qwI
2stByda0oSsAfJiLU5KeCE2r5GiwqNz94FsItoqLq+xxUHpmvq3o39q07srJtKz9bioTWF51RgyO
pwSmrg50LIqY6mBfHktCrk1gy2dkNPX2G+6O45QOKtVwzevHLAFT3epaEz9wUC4OD+xtKNgsttCm
g/MgS3ltJ4Kd8M5BoUjLO3VzAEDG4HxqCy0o7p8bOvn+6VTrjSg4L7KEL9OoxPxUEDD1LKMMx5hC
6mufKKvSz7DMmJo1yrQu4Avgb/s4Ph3KAIP5yJ1m9bZDeifAfvM/kpuFldgL3VEdS5adc2qTjGT7
Z8RcB4O1s2MCqRBJRTDPlQtmoHvS5+L5SUn6FUhlI9jzkxk3KPSMH3R91RkbY1AX4IEPAL64g8uK
P4Rw/NXzLL/xPdWitElPIyNCWCsZOtaHdEG72ruUl9uy3VZ3vEIafMTPELfrAM8zfJymjYyrvxYi
dwcJtP5OC6uA8WvZk8nFGXM9blQXg/yYBNh+ZTkQwLz3qzY2hT5wmfrAfNzBjD9UplTG61cV9uZ5
Qlu6NbvIumhtrXNc1U4uZklIw86Ge/nvMS+P8ZzTecwW6Q5W5pJosWTDG0nOb06z3SiBhsmp+mV4
9nMv0x23q+MgLNVW0K71EOakisPuaxtaLt7aiYlSyf4oQne9GKoCQk7ABIPJpFyGlZN0wITZeUZJ
8P1SFlt41rblHhkcwtSrffhoHk4L4e1OizYGoy0smlQDtGekIXqTF7OXfGEEYgXSF4nb7DT9AL+7
yH/LLWdK+/nJ0LzVDS3zggm6m7puSJlQN6eY3tft31mq0Y8CkU6lTbJH+UfniDMSRm4Jy1DSXv12
4UORHSJsbQYUGbQYVRE2bymwMhsktyQ7RV14ebHaFdcqQM8l/sRZ+t3Bqvs590NxXwXqFYuRZ5GM
sss+SPyeJMY6hsejPuo5TFSjvIQitAI4Nks+rb099w/HAJnDmxSvGsguA4UMSdEp0Fpiqy+7QAYB
ACkVOpM9gydwsXUiQoZ5qGxlgeFkfqsahCofpc1a4ZA5cBcPEDFcazHH2Z0ULNaqbygUq6gXMMTj
vyUJQTzYlfzAIlpjDPXkYySjATViURUvBISzip26GZkNAFWC7SujJIFczJLY2GZdJsZ0ZmWxiWUL
uNO2P+gOpNharpVuLv6CIXf+a+li+oKwGF5Lcj9hoTnJP4lpuOF0YbKyE5k+MIyhfILpSUr0jmqN
zCfiM2KGHxfoo9+8vjdqK/TwW+K26y/gs3kqPNMJfBLTCXjU3oM+q8WDeaZhFA7vp05XzQfAAGYT
gHifreldlj0FgAm3haSFjma51aFv8P/cVrMfsFXXWgKDUfpfA5A1MssZ7gkaaS6yEx0qKVYykPGT
DGwESPwOz+JxpwF4lo9r6HteDw1K/WVJmWqUtJbcs4Bn/V+bqLwfKb3cP5iTp/LtXcwEIqDQXOba
DrXTxc+iBlrtSGPFmPBqxmLm3pyH8vaDzOgIc1nfmfZOXXm02cjeYJmezBk3aeASY+YWT8HaR0TV
lq3z3cPdcR9wU5Y471Vt7aJ/+UN1DrnM5t/iLyq6h1i8eO6l9++/m7hYc7cVIfWad5lIuDFqZewq
YbMOiqtHTSaxDJvhGRyU6kl/cgMDFXCXN9Vt1SJVknSPnHpD/61v5PXbc8d00zDHu3AJookPaNSk
w0uoH9ubKi+qZJH6hfuc3ApeQ54Z/QHe68lMOzenCzM0QAFtL4X6LcOdrw/xBAonlc2jxMstO6zx
6FExn35kclejYi/XElCos6cIgR1dr+HdoG/AAiHBgfR7mVQuoXe8B0Xmcrpe9drDhucNXEor9gZ6
jipUjZvm1m98o0spueDODDe+FMZxpgd3M78nJ9V1Ey8BnIQB49hv16JbKyWb17STrND33f+wH2PI
lbMmEMoldemvoGSnoeHdbjR1jIDeYVl7w55ugL8kRcnV/BVtubjNPtn/oH8Rq8JSltpZoR9bbNvw
pjfB+z4qrmW4ZO+BkRt9dCg5Nqribh8fGgrrEew84CY9yiie+883eBe0SwgwEs7b2sFP6xVzKTdw
41iNr1JFLPBLTSsbpp37TMTQ6oRcxx+Lma1Xl2cNLAR7A8tM8oWKzvlI+GIqnK6hpsO0Vf/ZCCS7
thSt3HDhhetya93W7+l2xq0hQk0zeiarbb4Tro9EVJZakDBcZgjMaLF/K2v409OayHqdUvfQdhrI
3ALBEZ7juR4bHIPSlvVHtZHB9X+suF0YeQ1GfH3vO8OfcB6bZvfqd54ZJNvpEifQD/TutPjNd099
GxeOKCZ3gs/HKN1PgKBPApeYLOzbD5dmg7QvKd3rmMFomhO2Ag0Yf/Sd9RyXPcIEl6xuW+3t7AIE
hNCJggDx8vyDXXvMxtNQBRp9H6lqMZURoW5CXy9/EO/Xe7XvCba3nsHi3YIqFvTgyFlp3qN1917/
Ui4wRe1Q5LPRlJ7wd7trD0tSWtpf7Xr9CTaT8gRcL4JVHwRKKVzd64JfOWi6SQjQ57OHyywINoby
avHjkMbVGFI/ImLWXk2HwM4c+iBt8t9yIaFquS7MRV6cFNijuyuZe9AYs331AjFSQVMHveylEJY3
UtBhkyDkDdajG7yt6WutinZD8kgVJIIHHeUz8bTssSiOsgYaTmgjt7B66EFF2LOOwHffnT8tgp/E
TJTmBPMQTTepWEyToxAIU8MWM2cG0/I++grkn0MkZXZbvb4NMqYEIJafrCBkExFf/HciPNKSkJIT
R9HmEjI7aPw+Nr3CW7yw0ImF3ZbrZCTTGxtwrXt+JFrwNzQz6dwFa1eNEAtRJQPYsPULWK93WSHx
d8wQBzpkBo+aUKoCQBfrL/c/qXEfD3mR0VAvXwCZIYTLqt9uQwaCFPbhW0Q6D5BCyuPmL77FDwPj
y1Egjk8H4SuJXCMaTPfcwvqa/V/qHzPw5ih4Mo1onduWu5Ns+5CRuVCwPYfrf5+ViNhOFbGIOtw5
V93fklZUgl7vawb5rXmqdGNcD/knEa1SyBEKsUBJxTIsGYUaqQNbmTEd7+vj/b0a5BLtY1c0ktYi
pGSZuvUmAoUvngeiD2JcKUrs8U+7s/o3XfUwHq+mTGRLJq1I1kHq/80Z9pJa4L443ruhEO+CUcdL
YysqB+lb9dnr8/qY7qMvlT5nekH2lNT8f9ANunRvp1zBGLDNI4OUwKko0XlwJQ5p6J7yoCF5tBN+
dSQwB7BE3RSSDqyF/kD+kFVZQJSAh5tnrzKiBG1Gz6H+vKNohqRJVgVM8i12iE0inqioUhtYwxrB
NvfD+xRD5IrQmpd+Q8TKSJQrIYmjscgYIH7qVPX7HJQlkK8WWLriNFd+m8In4CcNq8QB/WkZdFVL
vkYRDIiKCmEI+5wqko2tG2NMQD9YnixcDD9E2c91r4MKssOLOh/aGhbgTBl7j5weU49dxV2cqwwp
COMLAzuIyzUbZ+AARcbcDHfaNdcXqDjdKpEOcC5cCUemg7Cx2c1TgFU37FkZhSuex2morhwr9JGV
n6uJh69G2sdUG/0BihZxr8TY0BIE1vDBzMprrDoOhT6/RC78qlH2/+oEIVZXxG+hL2UT2rK3JW6n
GEZOeJ3N0+mMarDlSuHXc0jE2dXttgPasCfnvS8b54tTwvQm0X1liG6xuQs+nMTfzNMyydFfDVNP
pgUZH77OcqFejTtK/0NaOMS0zGW7nHW82u/OTjounDFJBC3I7OR3V2zjbJtnTMDkFFyL+DvvzWVn
f9eZ9wynaDiWz5KUlDmv6IhAlHlN6I0XvhF67L9W+zUDbG3enbo1ecBtrspCRYe2BmlMUxWGWyld
6jMLUaIaWfMtPpxCVJG/HJZcUcHMHSb5f/r3Oc+Z6x7OH7ByXPt1A1Jiqg9TtlrFxlGVCVMUUtKA
L7q7pDUNO2+ak31Q9+h/2XkQ6R7wsnWGkdIpkf+flygRi5bf+Reb0l4qvMLRKSsvsYBpje0Px1Ij
dAkFiZk/LgAaNQfKCzn5A9gSGXil06DzgUb7LxT5EP7YhR/p3pDbfy6faJx/RsOzILikjAICtUBA
x/HEP8J5630RCsYU7R6FHfFVAzDUhWNQtf88E23uI9XXzGD5oK2KdqKlQToO8qfoJg0OB+sldA9Z
VRDFFnyMqhklE1+DTj5bPVbA3iMMMZ2J1FvDwBJMyKvyvAgi54iG+WKh0hL4JssjW1mDWn/n5M8X
kEAlGlANydiLsHqTJ98AGQX04bQ+DlYUm8npXuM4FuesULGSTTN/SFh4fKUYU5GdjUDm9xhGiSni
SRq9KeyBsaSATPvoEonysYoeBJO69NNUXxiANyV7kpAFuW3u+d0vTgakLr1qBZcUgcZ7juNgbrFl
EXYEIngcDyWD3QVw9cKmo0ctlokmemncn8okIpjBKfI3lAyFCuEHmGIopXOq5vQR1JRfDSK465mk
1t6+u78V140TJWvf95RKokbBXwT6+kO3xi/JWW1Ij1FDNF23YOrthTrwPxKf1XaMJxfLtSiPqPVl
gqomqAAvOjKq5czpUKqsxuwtxy4NMeQ9oS76IJQ7o6GGaC0L7w602fkhdaDDLkOmHLGZcmDSrUWo
dvSO9bniK38ZA83pdmZo+Ddv4Ya8SwvAkynoLBPVdnuzTLELOrHpfVk2oC2fvSpRSp/yVCPH3z5d
ZCYftfvUPPXgQFBItwnLRT9iI+nREyJqGZh5SRezDJy13YFqpJahBsxsH5ah7L8NkTSdwZh08VQS
DAw6Dw7NWHyBJ6ZG9ofAPLw0+kAcC3HxYWMe6BOsc+oQeqD9Ae1tF2QwmjhGyt66Hft83TBtQX/L
YZx+QbUbW2daUDzql6n7z9lj1xM+RYRQ0bmjdd4B7I3QVKITSc3HN7EDZ1+aQer4Tvf25ANPZG9h
H+0EAGwwDiTT6UpBPgrCHhlJobxop+13oWdP+zTfcBSEJenWmYQkKXp7lqilSrhJ/JKekKp6hDbL
wZWxrmO2Yc10F+sdoDh9QbzJptulvpcQYt2aTXMSMX/Et9rpn8g3x1EEP11fOX9PUJxc+ejUiVbA
q+i1OVT7/FHCD8x/KpeJnYyjKiASVy5/zDekbt3QM3Q0oNC6/IMrUhWUM5i9o8otoBDrIQsirOIY
64i3qYR6owPOYloLVk0fvMZ5ILh1u4sUlCqb29l2uWkx0rq2L7OgT/dgiGi9j619HKG+BFb/RLIz
5cR1tELuk/Y3A7vrV0rBkpV4FzoaKLSaZ57zHQ0itlAd6qh6XFtxzXpTl7qfjZ8wBFHWvb2E3uRJ
jEzvc/2lB1gIkkIKXTog2UQeDeZMUndiOwhre4rdwORwZaEiNX+PrcO325HmXE0R3ktFxT0YJiQ8
yDxN6XLsBROYTE0yEcWq9oxi4Ka2alNxDIiF3amu4ubTuGtOFCp9y3GXWbFmZwk60NxRGhdK/1aN
dubKnHfCAfcfcqvAckA4VHpuYpreTiJTd0x5X+bzpZY77ckXLat1FsJumwfjXbPq3qJSegJAjna5
Clf+oBCYVK+n8pmB5kX9YGJXm2Flgh3iZg635aiF6aLIaHyNABnBcVq8iU+4Qpfb1xx9j5dPOe1+
RXVAKnGNKbuQVxnQ6wd873czhLxVDtXf3Z2EmjZvBRS1zWpUQfqPtxKy2zF0sr1g+Ibzeir4Rfin
WzN2tDf7ruCYhwfGRAgxG10+4xl319OqrqxgkD01buYytrEk2yqOiriY9OBpjJPzldEha8d5/+ez
s+rcQI+bOjfKFKoM7qwGD5lVEm2mTe3ELY78cBYgvIhTRh4A4ZwzrWQAjcTiJIGRuG0U2Qng5T79
1lGIIJwLhgqspNVeRDx0YJnJc7o7xSpsIDhmJ3WGT8VbMvfMEKcJY+Nb3glK9g2t/8YAPLOVSEXp
gNkFRhOyRxFBEzzQsBdE928vIW/OdB5hybJMAmLojCjZjgRaITJuN574TjiQjvomG2K5aEALZrLB
jIkx+Tu+JbcTz+CWSj7883cf0/HYmH6SmiRRyBADOpwHtOAYgUAQ6njXRmRREqJ5i2/hhIbe9QEH
TfWDvfuy77wGGJKAvIy60EpepyrHXalt5c6gIz3N1vsP3g177vWvKnXu70YLHi7v9vexToG0mto9
mzebmohBI4RVkxjcVJb2UUIFCyJB+WAydc0232t11GLCu2VPHrBMApPAjcIRL299KRwQ4dY5bxeO
dTRyXoxPGWiIPTZbAAecRCuCZATvStvWOkDovNYvQGn60BZ0H6x5qj50eOwLl8v0g3rsBUmU5NtL
SG6SjIE14IZ+5PgiuiRTg3JOLrBmZaV6sV4O3ZJ0kUunPbLmzF3UeUMB+L+TSBi5YMo1IXbJc5xf
+tsBpJleYGsAAeWN3FxH20P7eXZlvb4vUY2/kR9Q+aCZSvdFVFBK9u4Le7dieVE9MJ/hZQcsIasX
EEpaNQ4qXGxZJPa7VSDSFB63K5w/8H+wT9tIA3v4bZyTny7Oo3DsYP0s92S177HlC7xOO8ZfzYpl
wjUzrA6bXaKmRlsJSH/FUJZnoOystpLuYaBCyUl4istjPW2NuVo9Y07+FDVKiHriJegsHBw35Z0l
eMA4QLSmd+f4GSdnXx4s3XjsXJoiGOYsIbdSNKHcmthTCBmZprm/9/5hTbB7uVzFujVhqcWcnU+K
xZE+8WMt8MGD8iZp79mQwez3znFnHJP5VCEu6gPoTREV8dfjTYyz3AgWle2rlw9GQb7T88e2udsk
EhRboGVeTeNi9CMpSOaJ3hqylFqZuC/nfXuD60M0d/CmNbvrK8sC7vB0OZyY1Q84fd5R1zikd+KB
384fHNtOOa+sxYecYBLAmQqQvs8G/h69qjtmK06lxYpi7hcVEU2ScB0wLvu1KEDBPsY9+sYVTwxD
1xW0zctAN0zephcWF+QpFChyYk9Yd8u0Z9W+fwAYcBbYgZRb9GUG2ItCd683P6TJrD9oYSakhm3X
DcBd3OIzoDiBZvqGx+Ygyd5fgiqJpypGXvJavEEv3IZ4VWJjTcasuewsTctOJpnKalb8aVy0yz0I
SAeLuCw46MeZ51jZ7VhhZKe+NKx0OaeW+uOhxBhmeyiRbDunXRRPdseVvvAOe3/IZwNXGr+kxxrN
F2srRqJnMC6TAefXGIZCsnR8mHXaK9cq3w+DGQywCgwm1ITr8x/qh3Czm7r1XXcpGDZWVT3jEC9C
0/nsORvTH/xaDSAF0n86g0FmshBPNulwze4lRQL24QhkPy0thC+zZl1pab9bl3kXVEv53Ev0Ongi
5vY7irrJIcH0jcatNAq9N0UV9ibjVttLmgy7ZZWMeFwWMQGlFNWcvhlYoJrjSMOt94+c1JAXH4/d
MYb8HMJXDmE+iKEYle3E3J1xPoQlzUjkeC+GaNpPYoeasEqk8JlKRNnxgx+6orinZWCSpF1S9Puz
5MAgbCcVKHyDj4Fgye/Wg08tAKCJkvcPmyxLwjO5mJcnEPa1NW3E7Dci2bMYdAj0p19SEtKYWGkB
uKnb2ieYrHuywA0RwY7oVhXL0WK0C1lK/eftxUZtrWYEnprmgVLc2+b/bqxR+DTiW7+4zfQL0z7l
Dt1Qo5AyhprodWBgX/A74b4zh+kARgcZD2qL2jKlFm/fdqiAKKD3Tqyukr9Klw230ohMfrRk3tBq
jcta+uzfSYgYOeX304HXxLxchRMqaL8UcPpGE7z3v+aQvvu6CeJA78Bx36dWSa1dO+oqMQ+4kjca
TrEm54MOzUL8rezaxfskIppf1oVrpJss3Tgk/IgmfyqAcgET1X+pl60Qm8mlWkWtPEWeW1PVi49B
V4Icw2R+UGods3abIPR+BKuzu4o5iyAQzHuX5lZabLQhGb+xz5jbsFHY7+XXJ0ySWWxAW1uipjUq
ynyTFZwGef+nyQka5djTxVRo0K1KiHNVGxbdRvAkQsHnTNycy9ND2j9x/URDi0zTIl3a1fj8BJbH
OUFLxk8OgGkVxftIm6Dl6meVCG+qTMJrcXuW4/iVWt/hWjoFuLSXEagS6yfBAbP00Uu0/PVOFHfi
XhOFyY1NRryhwW1IoIjfbQS3ttGJnT9OWeKBpupXC5TQ5AwnDjw6JPFRemPQPIw6cGzm2ekjJ9D+
LghnakHbJV5xZDnHF3is58iuMwfhgi544l3rHoMT9enAkFhmka54Dcqrqg1CryxHHC/M9YZoWBCf
qZyxD5c4UmB6r9UNHeg8YRCkShAPW6d+GMJI50ZYVmPBnQRNceyk4u64QTbUcbyh5dLo/JTWFpgQ
dLXOCgr+m0OvMSdYJp2oeuo5NElMX3WAAVezFksT3/7g2W4KrOMRk6zmWrRCsFQwon945qvhaa9s
4+50bormPp7zvR8RJUq/pi9PgOx8/gEJwQuhIBx8I3ciCpTBNI3REWS5NkwqLG8s0L9NEapqTe1r
wkvmmQ0Byg3nSscW7hc8oQFXSaTihPkhVTKlMW/e8Ud8YJ0RCrzFYTrFp/eN+aFrK3N5GsPqZxZa
75W7Tp9L5EfsxmpOIU7PqW5YFizaXKFGI2KtNRnPxnNhMh6DMs7TQLIfSCqAP0kPonJK+pHm+3EP
0ZFcmyw8PoOuKLsCKS2m6kJ90vcdCQuYw78i/ci/zvLoAaMRqY3wPwUR6JHZ3HtODPCaH5OcLSkW
wi80zF4NKdmsEIdG5cXsGGJPC3dIZiD16KEwZflMcWDxV8kjA4x0spIx2XpFXoflxqpHfIxdrl0X
ZZqFSMgVkzwtSrYQlzVKUSgJHkRhGSOgsgXBKJwrhLrUkgL02zYv9FaqBkMIBv4vOasxwdSpemCs
zuf6b0YW+Urn+dTcL3NPCi7oGIXp6dpGDF1bA/z5qyVEpCV0lyHcAdQHITKt12dF2j1k2YUVAvJ6
rbCGcO6nOxLVifc0LYDLF2NpjcwlkF/6RznzLAIvUABKg6YAYHsbURCMsmtEjv8llUonYGPQY7Gu
UnOChWOUv8S/OZAHLfcrYlx6BulR7LVDeY7L+0uxc0I3agLY4jDR3D7XsHvuB8iO5zTuHzAiVVGm
PidXwBH20yRExX0lNMm7VCpXHMg86iTqOS0k+p7MTzTNWOoNCwYlwCTtwKaxOpBNCDOeSfkabHTb
MGf5A+Yzr5SOll56ESHXxtGH0sBG6HCAfnKD4R8zLwCOfpTfEEdQgvI71NGbxwwzVxxSVwiFqqYT
j+mxGMpYiX0zo0lhdUnPpE8/GrCsiENeb8pSEfX9yW2G0nXmWVLOREls7s7WCoqQ7QiA88O2ZfV2
lk63rW/wGdI8hateAIHAU7dzeJ5DbubstkMjpAULSHNuLylvFGwIlnjJjMLD/j606L5l/v6JNnth
tD3ngNghzOceV7bSVILXNKh+qwieErgpDAH0fkXbDipQzI4uvKGaXypa3fBkm9otHeYGLjE+ELzk
6HMVvu0b8Hbiykbw3DAB46bT/5AadGFRD053rpGrHfRH1f8cZwa+qtQa3i9UVVJp/UfiWsK+I5SL
p4qkhG4XkYmfnJ2Y2CKFkgiFqY4v/l3LQ7CPzE92PBIMzmq8vF1iRrU1O67mWkKjfTTysFwBATZR
im9xL/bPXHeMmHLpgQFvG+rt8ojT0qT2T69pQcXKdwPzxbr7NFR3xxgsQ2QEWZtitr5OKmdrcPN5
xmhPAWYP64zwTt9NAFPTIW2k3GUcQpFnLyiNkSnrbqgnmMxLFAld9jfc755UBX3SFAxlQbAIQSW0
bj7qS8d26R0RzfjJczsol+D3sn8FHvkrD+ajQD5pUAISfLe7lhxvlgHrvTRG7qo1bi4g9ZMM5wBF
z6UJqg4g3lRTNHnK7vNYpD+d8HF0RHFNaLfRaG6jiSlWrwap4Vas8s5qnhvoWjhQJhfeh6c3U9e2
1Sj4YKO5IbyAHJUPb70T0p9mLmZW8b67yIDLuJ3p9e85ncRkITnmJ01c4zKclJ+cQNX3zDQkk6Wt
OEGduuPuCCrLo0+B/w7GIJPdEy0+/+uMfhFWDCdfnIgfLpGl1bigKID+A4Tob+LH9LFwplNpqbLK
a4IzeQT3OSR10Rh5bE79YWwaaCLmD0IACnEjG5NLLpnrCRVxrzn/S7EfbbzmzXMSnjWAPHPS8qih
UvyKFg03sZdRW0R0Lnqjxpi30JnyqpBoCuhzmlpQUjFyy0Cs/BYXeWt/Q0cpep+vn6w3spUdnQ4E
uLyKcelwnrpGwbSn74n2amSb+Ou84pVrQXDjCTR+KBbqWXUipd/bDLBFgHQnlPaxGoi1TzMHyeYt
iwHh6Tb0ZbyhxBJFvjr4WxXfZeCe3sQX66tjrJ7FVTzFxr4/e0eMEqijnmTiZ1un4KDPaG+EY6Lt
Io9gCUCbFXsw3yGODtA7SYtSsGxfy5+UKgH9f0wwrEKYobNg27NAIavMoS3BrFZffO7+m2rQx4n5
D9eg68AuvCHCyKAd+12I3+uA4s+V5rgG1dVVb3+Jfuu5hJRGo1b5NzGgSJZEDHVT9CRgCpr+rZ43
8Iu+RIUOiXnvUphE3+bbVywzOkAO9CeXMzuXXuT4MOODxsp02VAbOO/ddePmlPGPAGx4IHQMsbR3
lBO6xJ3duNBL9LTa14ydAu3iGYOMpVHC0HkoADtMSVfFaZPwDw7n14SXj9H29FoCWBpIY1Iwb7gl
zGzAVB9ZxuAv1W24nWu8vXV4vCqFi+TvQnYh4LZ8VC507ND2muOz/bngR+K8LhHPqxNGT9+PjCk/
ms1HdkVO7CP7HiRghpfHBDDce06Nh8/baW0E5W8bh4xubRoDkWwexvpdCfKPqDTjQSNTCvYxhg+r
TrX3yNWabGnMWudPy+jeUxjDeenkp5/uHfJ37Kf4HylRwJkxMONHgYaQAeexv8UIJy7wc8K+HxTi
gFy9YZzYcuIT8Xt1xtMyPztnADJAT8TdalN+ZdNpfQKYKvl+yf0Wp9m1HlHvstUDhUMJXcsVAXhO
uO8X0zAVpiqO/swQAmQBQfnU2Ih9xZqcotKUyg15/q6iPLFNj/i7nL3e4nFm/UgRrPXM2ZJF6GMF
9eFVHIfGurhHsqdrwyiC+uCiHW4B4ppnuBYfjiBkvKwSUzAP87dbJ+nhuWQSutJQY47C98T2Cy3v
84sv6lPFOPY/lZlnMtWwDFdFMOwd+3O3Uum3gUirJ8cIKEBjgT8gYc5U4A6Oa7u1a4L6gQykZiqf
+1Y0Uf8ZvmDuvojnOiU4bDJZlniFK8FaW73OMAthQ8xuWF0ULy8fGg4p65JIokIpHUfL+KaaX9cH
UUYeP9V6EdzksgMJARkWOib5YcDvStJdOfi65ZoMLNMsOMxxQ0yVoztnZatoIFd05EhgwPsB7WjR
6lVjbpxTGKWwtfGC7vvLICN1p812UsT2HG9vcwzfGTRBbi0WqKNOy3d0AkUUWXw2UH/A46IquiQi
Tc4XTi1tJBSiIdkJjP9VBxKqs9SAWlgLDEC+pfXwVp/JzH0nzg7zL6CWKSRnzJlPHSf6Rir1khwb
oyeevnb0LxYOeHY06JLk1MoBJK9WQlogh7Ad52qzBytSg5DtZODUIdvuztiCujrb5hngePUZHyGF
R5Xbmv9l+dQYB42bZMjTSSU2JSAvnoMwgsitx6aVTcGVtX6bQiYVxhiXC5IxF3UwVU91VtP/iRrb
pup6j7Ko1GS+TDxiB9jVYk47wl3agpBVkq5LqzqBd0ye6Jc+fCLCQdt+CvmgvSoL29CdZ2DMI7ZZ
YmWQchNjFVTLCxdjIH+SIDS09H1C+vZCM874KNz7Z2/60vhml9KxfVAREvLEJOf/+4sck+w+l1DY
w7kLjquKQku6aToaFSQVFdIXfy9MZ6ncp8p36BULIY7vDem/qYdpenoShdumEt5u7htbU6X2P5eb
dGhn/PEGr2Xx+wsvFo6Je5pI+fyG8cmHdD2QTnU8GMEaRj0CwkU7l5ImwW3DT6DBUBUYDlyTmmC7
qAN5DnFWM/fdj1TH/2ciLx1gG1YnPQErcSUkEOno30J6sO3ohqe4/8gxSzsJqcvXg21RTZFGh8v2
Cplcxhh17NIxDPyxjJO9rluEkCNqWuaNs1cF+MHikf6X1M9RNwJBVWv+OBLZhV0h2wv9MMH+Icmw
Gstt1sU6yy4dWsr2oO7/QUjRcFU5TbMmCgKG66AVVGSm8ylQ+Jz+nVK+N/+GnzXMFDC8j7rin1Az
NxTBWkg51zVrsx5aTgo+/aaAjkB/Jql9KQ3GTT3nbp7IbpLrxBWcG8UPMu0u256mT+Id69F88i2w
2LzhipoI4kouyHIGt2uxqP7uyimge5mpxXpyMYK32iYeum4dmEZ239sA0UdKDnMtDxDVfzOS74xH
xZOireQWKZz9SwYgU15CtExAwGrCVU78KaCnm/z3OX8HUH3Dm4cNFUEsuDXidWf9MpAUz7bpFptJ
UndUWKkGdfI9XRTLyfu3gKLHCbW/9TKgg/IBCJuyYDLPqoBOTzqI0MPg+tQFQ5L89Zq+1g2jcDg7
5mbEIZapx/c9QkV6fsi1DpC+X0oZlwGi8FKcKvqpEljgudwW7Ma/TRyX4Gdk0lcWmBFzjoZQQ+w4
Wny5AC2omc9XY0jv5S4whEzvC4SHqVQ/uDuhlfOociV/Bh55Pd/43iVL+OtSpQn7em4Fxe8nVmr2
F2FMZY7xaPm5mD2FJswTFwswcTsLS8EXJf+BzvBhIWHyf64uQ9D0kLkLPj+9hdiDjeNXlFRCaOBQ
eMFPn/tdMFOuLGC66WCB4BJRnyu8xe4HRzYHjor7BeRj+/uaGZ0XGB6JxMmSqifdJC6w9fbUxCzb
nrt9Xi4jCi9RkREdb4PK2+NfC4GEESraRKwrCF6ypIYnrbuIQoN/fIjvjI2xhxgrK24Ssi9E+oxK
XAm5vLtzQFZMcnffweivmzBDKibJ4EjfGaLv/J6XaFBG1O6qLVZRN1oo3jXFJJy1bzU0vZRbwYrF
vuwVbXuAIeQorrLwGEjdbGRw1Aohu/K5OhB6UuI8xM/DTnPLzd9uzQ/znWmZNiY/CXN3a2Xv7RwA
KWUtTLtVjZFm4rE5YjISxjMSQpzzviot+1+WbzpBHLirT4qbKzyAfF4FCzFao5l9kdUwYfrGSpiC
WI8+y19GpeiiVxNZtxbVRAeFQBlxUUPKlpWTiCdws4egiCTsHNnrM+73YN/Fr0ASk++hnRss7yww
SZBPdQw4QyFKiadkiZnNYwroBYLNVg/fC4vNQsVRmq3NQZvEgyYhRHuTEN9bC//Ttk3Ii6o5og3t
hSg+0qlvNN3e/oyL8d4DHpcfvLGaggR40yRiGFoQ2ijsRE10SOK4zY0XWz1c2Ul5T/qcq1PjURSO
ShJHhVlieWEnJqTIK3+NmrIziyN09GVASM8MKJIAbYJukSvMoWZQtvA4BVTE9yx/PJJTOx/2w1z7
9GES80guZHuWfOl5522D9CNyiSp2DC0UrfIvhMjok7gYIjoPvOaLm21UNNykPVVfTgpANjh/e2OJ
w6VZkEOMqvv8E92Fj4VseDHfQ+6wGqvmKhgVyUSln6ikTHVAOXKGzrYJAvKM3BOVK4dCZNzqT2/Z
AQzYt2TSgjhJxvmOJGVC5lEmOq3Riz4J0T3oKfLUMApG8n9jSs7c1zAIzzGB74lMQao4F3IanQJu
F9c7YWVYLTB0S+3GdPwJ012oj8azidGj/UCZufdSbKVk4imZjolS84pJBPqWZxswCtTm+c1nZxld
cjBTE9dDkf5OmwQyT2EAb+g65hJe7WCsrLzOUuYHNCMvA9w9o6GPE2TVIXBYwU0dBeTJaN4UKUSl
P8+iGheqDIB4znAD+WDw+NpGgWzWIttyK33smAkG6i3QuX8Fm0nK6CqbxvfGHqZ0RPpeCrcphdgl
CUtikQwaivfnjJwtH5dukCNPHYw6Btc1XT8W0wMHi0KMIOw3KQWnVV5WcXGWpu4cvpzqiUhDMdey
rC9BegSl71+gLTI6nUZWoTkGd+1I398GSUBCasXmk3Gr5stdk0vFC4rpQ8uqmnQyE1qoGnDrh/iL
w0dr1G/tQAkuMmdbsWimKrcpb+/3sdKlFHYAnKvGWDRBzvO/L48rix8vD6VRUuHFIgz4awYce4K9
D8cg9Qu2XLRD8ELOahQugR8h5e3berJGr/8sEJBremQKnvqbCyGA9Xe0xEf0z7ESVpNNeHmcRbeB
GjlYvqpHzE3CjklkIV7msalaZZCzMPf2pC/p8+5cxOYrC5GoafdIbYFtA1SV/88qyAqU00polSIX
iYVXyhbX3VbJGkN1Pu2hogv+KnAXwfchjCbJPHBNtDQNNQQQXPElZmDzJtzfdy8GvvYHKWSwDBxo
43pA9NRYhJiU29FSkMIVJ1Kn3M0Fzd6QeTaqeKhDVlzT15trL/kGsBby+YBGYu5rXrDyxIg9v9V3
LBxk/iGbI5m/c02d8dcvP1tFM5OfMB33DK3wxxI8OCr3yl6t4GBXijKPC3YJ/0LDz6YwpwnOjnc2
oIkBWPDHnmt2FS+zCe1X4uRebxIrT6DtcFFqk5AH93BRZYqtHkmetv0QocLQ0SJ5c+XDP0w+MogT
CHReaeWsl/HPSjS+cYPBqUdEim24Kl9jpB5mbaFxdMYjfdEqlm8IvpUcgQU/EzQq/GwxC3HhkvfJ
VYueLebw/xA+6HzQfULAQTQ6ChOSDnKjLjBb7ZRytf15AKsoShILt14wFwzrQVQdKkwc6XM3LLfK
cSb83JeNK23NyIHCrY/gQ73xUkv2l9z0UmJBvP/mCpHaCCAFJNOoamY6ly36zeC33tsCi3ezbQxD
ppS8oiKV9uGPVQ2oBa/8gJ2mYtbJ3I9T5D2nGfdk8VJUcMSOLOzdbLwwvd74pVhCdMogpx4DwCDy
hR2GZbiQmtulomlQN0gvy7KZKxcf6/dtT8JBmLxFOn/FHIARM/TMFT4ycvxoSvXvIhUErXxKSxBU
JBAw3WzcXewDWlUxYYO0G3qJ4AFUnvc1ZDvQiEPpLFtA/P+yuVIu9cQI6uzJmW2Up/uyQkIDHyyz
gANshzIYBW/D88wPXMHOEgigZC1Tqbv2fjhrHZ3EZtlGwT1mWkzl9oaSoSI4tllNnUeiWKacgDOv
2x16jsB9R9v0YDpaa9/lrkoqX9osZE0mG/5OtQ4nStr1PkRAo0KtiOUkINP1OCKUNHrzKq17OfDV
CBJSX7DrxHHmyBa0touJBrzc+4MPR24tU+LakOzAneU3iG0S98fhaRsXKbQwr+QRvHCn74pJndKK
D+k2oRDLXFOe/DtTAKty5G18QP6rtXMfW0lsQjuppyeGWBstG8UQW2Zf2txGLw4ysGE2YYG/XP3d
zEDn+NpmkTwsLPj3lzX9eWRDal0p7xbHSkZnOTlTJuxLWlUV/bt06OAwLrNJmtgErY5XAvG8cBwi
toj3xtceNbLbMldaXnS3y4RbnEUbArjxcy3FfdW+Vxz1S45GV1svZ19XverbHQlAzGy6NDvtSmEj
00hFfEVOOWjO2JcmH7pFPWTPwSfi9O5FAfp0npQKW/s7EzZLE1wnv6ULJL7pCL2Ygv+LnTtIXlsj
dgzbZC9A5kNcvuVBCTdHPnvd2pacxHjvitzHDkQZhB1lLggr4pIkPhJvPTvFwd1XFZg592+5UFQd
sheVMxj0c7hUi5d1o1gK5LsU53L9OfDZ4EtYN7yFwwG7mnLeRzsLMG4A9Ubvu/i53nwUA1J7UB0i
+8wpajHsW0TCkJeowc739Bhn0irngHPz3Ntl2Z19A2rxeQusKSKFlDW2i5gYwvAqhjLp22fPVS6u
GDUN0B1AWutcH6oxPKPOROiOx9LAlt53x2VqODFVv4qjCMPeWw1kt14N7TFppuYUGhFlck9IFJWk
5Wqf1vxOP3IKAv4VDceYdXD8TcvEqRGTu+4hqna8duhYfyKN7eZY8LGzB8SbQ0wy7KJ6d5IcFYt0
gikWG4YpwxxPBTAs6mHnwIsGSDpPz0NK4fad+7zkg3PrGQveTwmCkEHC4wLuxAyiU82GMTcxnR0S
YXIvBxN9qUDpRprrwPFVnuH9HfhQe5z2OkfdtPyuPeM8mjeFAVzcFq2GYv/9cfuWddmsKYl03caj
UBYSLD1RpQ6Zgje9nfk0Yr2Maq3yfBaj1cGEbzfdiAUxW7zNQkEqWdE7bov+wqtgSoKghNGnMIYC
wY1aL3LJD1VbZ79Goz3TJnT30Ln4HoVC/wbLiyOPYJIVg1WPG7zn+7x1E4xgU/l/1Rv0ygRQnI70
3KX9zzzEKYa4rXR4Ag2s5bzWiHkwXdGSbgkMXHS/O0AKmY3O7dqk3Jd3zwrAABoyL/TwDZE4s2kb
aDj7iJ0t3xNTEwNAUOTCJyaP4Rx1K8QyNr2VTXKDCmbYaN1VhdFF48CfbDQ/l754BJxAJRPuAiMd
FFOZJsAfV1TpCjhIzF4AlM0yW8HagyYSj/Ov+V4ar+MIQX6YqC5dVMRtZfckAuyvSjrUcrbdvvm+
R1gbF/+tKE01iaAtoXF4vpzYqSOGii2Yc5b+Vsp9Z4Hy5iEUagZYrkq/Xjh5iBvxtvQwhQTTv7MS
t/tgCGJSD5fedH0bjuNW3zCdhC09enHwum2SSFa0k2hagMaBkaONKcGcfhqAr8aFXcCfgl6Y4PAL
BFA3T3YReY+T8MKnF6f8TTPRbZtNQyVMkkBA+fm8mbDyNh3y2fzkhAsTSc5TCZTH7MDWp1qnL4Qk
VomQQPnMFJz+ow0e3TR1vEfw8U2iqGtXQvwxQOUXaMibw7jOsCuPIgT80PNEDH8qHNbm4jDnLyM2
0WHbAeoXAkUvLOj5Xq57ojklXoLejEK+f9/ted7ZmEKtkPbUBr91i/OYKNfFr3Oll42LoQV/rgCs
YW4NjVWCatxvUOx4FiwN5+Pt79OgeMOLSXmnvm7MGv+T1h7hHPWxibCT4W6W22DXBu79kHVplZBI
OW/s4y3XOdBhsbt2NED4Y+jmN4eldhhgMV0ibthraI7X5UzaorRiqZfzVcW4smY6M8pAGp5X+c0Q
F/fgxEot+uLpm1hY/o/HxcPAd92jcQlsmTN28iIb+chdnN98xjN8KihbgCI3yBZwlQ3p9KPU4nXj
/ryZEk04HPdhjRq+5l8cxnXpR/ueBlAiQY1jcE0xjB7lTFa4f8AQKo6XgJ8IGSNDVZk/BM2hQAsP
ehpeFkB8+Z8n6I1rDLxPbvURWJnGv8w5vt7XBy4/fg+plFfvJtZIOTrQFaUASSrWFxmyYpAwsEn9
6zFJOKdNPnc+0y5R7DoYmAOABaK2CGP4Vx4jLeTOqybQWFfPVh+QX/YYb9jgoVSZkUsg8aPkx4sB
kuQef70BJLhr9Y+dIkdp91Rmelakq6ZmzqbZ+bO2COavmOe+aPpGGKijf7ZSicBeW/EHyXAI66q+
iGJC6DzWRKWSEKZ79t2c+mz/qHotu9tHKfk1HnEYeQdXVHwzvWruut+Gi3pfmT3Ur/UUaumtPBXp
HR2FFUp74zUOwmjRIkdFZwXABAKKsdgdrcqC9BV7qVF6csWtJH7dC+F1gqFPjVXUD99aBpkc+2QO
1sKsLDhqytlokyfwBaW8/3/98Brj2Ei6hTnR00l+PpP7agLI/mP/gRy14+g4Ev6lrPYNUk7tq2C5
V5wsCMQWb7nHvWraET0Oe6+khXVgQfQGMQDq1BtkfvIJOU/owByH9u9b/0v4If4CeMeYM6SCGRRX
PpNcMu6BvlKaSHvsQDxf6wcLjXEnq8lEhQznff6sFf9wNggLas98ZoZazUvVsTT6ciXuu5nIok5z
izM/8PcCYwteOvxWKPFqwzcj9aG8zLC+aJJ7PaHD17A7EKN31WgJuIv9Azn3Xoq+y/2nqY7Nrdwt
/Fyg3oxsWqrz0EZM9w/QmcVrLUfMrEkN4XoKhBM+fFdqWKM5zE+25164XMJ6Z1AVcGGLX0K4/SxL
D4bXUCuZMpxjsCut9YV/eA5zWYPntrtY1Dvg55fhuMi5sIhOGo6G0mK5laL4ktSD9q0dENviW6zw
jAlzX3hq9xqCKubV7ubh1WWh4NG6Zk4Bx1WAlUKyeB02dxlCE3zwtvTvR9z60NsdC8WP6kTy+TfY
/Mlmu/ZVK/b50W8tiMMsUa8F+pnfteKav2iCDJzzo6ZU6/+o6+79V1JaATSPZ3ZsJfZ497O7SU/L
NKOMBAr1LRk4lrL8dU2NkD1eHUvwLxc88SjYD7iWRMevWIYpeozrifdTxmesq9U7jTAuvUQjsvrh
MrpCkjmreoksCE324IfgXJuxvPHoDTf/+dqGjW1yTDujjY1Qmy5hrcBDwxtv13QVfHI3AtbyAww2
zdyu2cNG/PvmRamhFJZ5h30zTmiV0SfnHuM5VV8RG1ALg/lbP9Q5p7GfpgEHRzTBiADShT1eLp5h
KyZDJXEHca8fjcBbDKb77X/lF+czq+AFHQJohK/wMw7hNvCYTFiKuCYuR8z2ZpaqaenMhBQ0Yc56
KIeVtW/AdawSYsMs5UNHF9KHdpjFmW52+O0rtQBl0Xy3jFe+fc8+zVQREszzZ1ETprRYM0+s/eos
1PdClw8MBbEdRG5kqwvkdCSALLqrdZV4JwJVbf7ATgTnsdZ4g5+afV1+t4nMkAtwYKEQcxkZeQxg
ppD/H6MvgbDyUGM1dCqowqevuOTFt0aOIkGv8PmOr66HcKrrg5+7lLJ1MNGG6e620Jqhe0/Gc+76
siqWN66wj2vkC9LBZXbghF0k9V8TVdC5pKWQHXnMJpZf/xs+xSWjDndxckm/fhWQaUXslPbRg9wT
ZWsJTt/jXTicSA27WZuLrQeT1g0qBYh2q1mcZ8yGgQ506Qqw5Klg1tcfQq86urcjkU5oBtHT3n9U
rBQw6Vt6xHOaB4M0VeVDmf3F8Fh1vDKwPRb8jwa0KKJRmGNCqQa3Dnf7c/DatJ+8Z3j3EuZmYe8v
0jCt3OemZLsZYMRuCfP03LvwVotzg7OIc2G/cUeP2mw5H2Hrq+bjPDbvvn0Nqkk6tk1U6dwWLhQO
fhKxssig2AIoDU5aODmIILr++ulk9BEHucf12kYj7V7YA8GyK3WvrYRvJwABx8ii7FiCMqoIE/9a
zNMfMMeX5RUGj89D2WwnCveHbjrUyn+zJCT49YF1mEiA4h+vBif5FG4jWvmvJjr2QDTkXsMykpu3
Gl/soqPRUgXzpQguD2DRky9gW0igZSRSDXmsDCD7bMBnknoRwlR7lk7Xy7kI4t+wBPQa1mh0cizw
/vnHZkSsJBVrmQdpLxQ0tg6HuzvgVsdj1mQGab31xb6j9NE0p5QfLJUREVeNdzzSWgiqKBHN9ID1
80sZqVw/BSSb3cRJHddjpuCuZLMBFbegdJPrFPgUayQsoYBfdaDSo4e+u4TzPO3dDE9Thl0YMDmk
G1LBdvS5lWuDizlClTWdMqJVUMvs6dWzjtrOwDlsjyja6JowOYDeM077MJFYb+ZslYs/KI7OW1Gs
cECV4bYPD3MvtoIv9NOA+MR72as4a6DMyf1iVkyv55RXoyzFeCwOphmFHfcx+fsRx8oMmrvCyxK7
QNbLTEN2MIz8B3J6Phg7ZN7zyv2l4W5iqv4acgfVO8LBCSU62ySUmLyDaE3kT92LuINn+bGYmj48
vmKR20fdAgZsFG/s3MUxicE20rVmtsFUEo60Hp1nH5eTfej2wdWs6cflv0ookLPzZFTDt2h0z2ZU
VQSODzciXHR1m712gaRX9Rw9aEIlM60k6V+vHudqgZwzTbDTbE8e+8rQ2svFs77JrN5dAZ8Mh+Qe
64+N9hmUYc/pVl4lpe9brIHZI8G49hLGmdZmg549PYp9zMiNB89+BIRRsSEwedSstQM2uwyct1RY
1bLxrPj4dcVboF/ut2KIt2oSCu1ATWsSdxdIKky+tC6kSb3bzTk9TpzRMNl/koxwRV2YaHYlCIr0
Fh5JB4sM1km/rJGyOi9i+ZIBFK28LF1Zk+58VLN8rYb1uJs9v92rzysVZaqwk/hfuX+K2hdKNJ/A
l02hxUL/P7iW1gN1Uflgo4ATkEEYqlM9r0s7gO0IEBenEDtNonKknAiYG0kOxRn1YJibI1lMj4Ud
PW/OrIxKs/VIO2eM8NaxTisTaa9sx85kkTLr9FuqeXqbNHbFW06qu88rj/FVSIa7Eu09ACAtiYBu
Oan3WVLRwlk4pMy5nezRX2e4CYpMSgJ56uBVZntzOpMulxQ3T9OCGGIDkf9yY0POFxTu3oVx3LKM
ejFZg+nlTyzH8bGN2GqqgFDRRv62tmzyMjzlpPO3+E99nFzcTIekEN3B78kwh1IU1EXk35MSy0AD
1BexI4mmo9Ryl07WI0evuPHT+i1RkzaIbgrVG0E0YS1C8YOTIB5L7H4KXWPVWpIadOAtkrCazeDJ
kB91r05lF1IDEC8PbGGuv6mt8WSloAnwMBNDHQqUJeto1yFrsOrJpYpesP6P3KJW8Gzr87xzV3+R
LSrVpELnv0I41XuDJIHs/eFCmTXhdPnAIgosmQgBdog02sgFZ5mFRmy63avujSUqxhueAp4nNFoZ
9IgJGQPyFi7uvyZkVas3ddo3lEwm4PRkXJK46035a+PMFsP10O86pNGvTa8XJHqGDMXWW0G4B1Ie
EzsHNGUGhaCcM9aeCMvdaONTuUAE0C5/jA1EH1dCj73VGl5LcMkdoPJNArzrcOOKLe95ooxpYJBu
www/SI4kNz2Wsa+0nri5cqeMGYn470jbm/k9xe00BWf+HU2Hm2FIVt9jGNLJia/tSQIa+pFhwZYg
swCdfpslhanye86b0BNoPMU9nBlTYWJyhIa+LO1ZEskvo1Q/1zJtFb2m1bCIN4QatfF9i7AICLYM
WNhzBRzJ20zbdyny0W1CUi/2H1tdfSopqfSkHwzz0cuecn6DLWXGccULsmYqBPBPwO1KP5IsvuzA
b0zpmsSXStZLQPX1R3O3KeZcE69o4u0ztgdBchIPxXWD+N0rg2EP2+G93myABBY9ljXNCULLcMTY
yIXol1QACM+bDp4FCRAgLPlEiKWX8kF/3v2152Uplh14zNkgLujDcME6tMkEyrPKxGzb86TkOLtq
yJfjIellRA6r/3keXLQlTc3E0CP4YhMQlQ85mQnl3QohYIqf7CgvBMj9IfUpTr73132rzOcwyFct
zV/Ip0VjfiJJwHR9GDQGlUmCEcQ4Qgb8ngu7R/MyGWMWF/spG07K6Dll3MufNTM9azw6s56vQfz3
CS1bLbnAvlvFnYZob9gtXOOjrbsf0iyWOgWKa0KmwJ5kmadu6mfyqbgLRXLCpTLCZibHW1h4eLlk
cPtagk/DrMdKI8+2brYWQT8rtfsGJI8vde94WgLnkLTibte+URZFy7koaXucAc8f8Tf8K4ilWGH4
CcW8yQq4eUz4z180Yh623wstkd7twfZMY59LXa4c2tQVQCXpJZbf3FNTCL+iI5rdxoSyCTL+RlEp
Zbt9av7dDThwpp+HPnOEhFa+Ly6Wnuh7gBKYB9dRspgFL3r0BgN+RNGV4+hHmUiACNRDxvqdzBmC
uM2vI4+VW1i8GsY1TRtEVhEoFQzHRn5mIiqs8pgjlrWystncaDdSXjQNj91/4yZvljv0azlSFq5T
3JfZyonys1ZIRJsmCMECWGzaihvrTPomzEB5AA0Vba9UjrOsVYnsXXtXyp82UU13z7tvHtLD7oAd
KLnWwCLEMRR+5F1yOIZOafawJuzk9buFhF2xcK1eLHmLyQE817/8HTPWhmAE5DfD9zYs5dqGD9Jn
xaTqoTJo8qvj+wOr7fsk4Z8hUoQqU53FDNh90gSKXEB4p6XUdNJmqGTz8DU7tLi3U2LXl2DpLJlg
mrMzXteAxdw9FaQVnXcJrbcvsU5ampSXMqm8fVC4lKbfiQSCEKWOSilkgwMhokWC9tTPnzRsy1oP
0oSw7RJzftGZGiMP1uD0GPRlWVRiFfoPNJcep0egiVp6g07FtczWpsz3CuMiCF/lz741CgagnNY5
xraJCiIwndk6Gco03v8QJYLmNcBguaz5o+BRYFioGZSrH7S7BJfNeHjJBVTx4GjCLJ4POjRIaWLL
koArO8haFnLtev16yBZbHIwa94I3J1GeRz1k/FsTrrz84iGTtpvOSLnwBhYd7o1g8b29XVn8aFE0
7CljhveMBJLbwQzowcUt8mAUtuPqv9b4rjn1EEdI4gz9soeS72Se1PYHqACnA/paE7SwTzI8C7gN
a00ShluhWL7sgjAfdKQ9oA6FCXxRrq4+h89rxl55tYzQCN6fD4ISgCsIE4AoxwpxtHIBgN5+5uy4
bnvKmQm1Pmf3b91TrtS52LZh5LXhbCGgBr7Fw+9AtsnPgawRiQRBEyYb6ysyWI72H5CUspYpP1nq
o6lSmPUoaCdg+D//7dIrMoArGT0mm0afUQ0oMGLuo6IVCDl7Dy4BM/xlYj0AxFyW0OmL47Lvrawr
olYbh6y7ZvZj0noTcmORw/g9L/v06Z/FvZJhArwo7ji25Ruk47QN/J46bUH71whjEB4MKH0rRPvB
d4bTYbzQ+AjMZmJynhhLQ1pDbIMCUD6/rSeqsc35JFFKjwk2DuRDM2xtQhGCYd0hDhlPzmMjmt1B
lzX2WbsxDnZtQvdmTwTW7YL67bFZuEg4KOUYijAqSBfoeoHNDpzDHD6jksdGmZ6TzufhI6+YYCRB
zB2C+vCIvNb9+mreKom7lUceJ8WLMm59oEDLzSjU1dnP6T6rixcioaCEgMXKRJehKKaUxkhzWy4b
siBw07Z6E41H3tiJc4OdueEr8FdhrK80WyWlsoq4GbQg1lIG21hy28+U/zTC+asMo5pe8tm0/aXc
xq/yK93YN5RIrfHU/5ODZEbr/0Z1PwYcVOwe3XITzwSwc1wdFcsKVaERvKFM9ofhlc4vm7KZ1GRN
nerO5vUPQKgnp8z+HcoopkMyuhQ7a5iEb+GTXeuw2tL0rvrH3+HtzCQ/8ADJ33Y9ZjTdHEo8hstO
84lS5ElywYi2jk+htDQVtzQsL6Ey2luwGDfJjuuAQ147aXyHqwX2r/ofX/1hxnNAI+IIYE89dtNb
qDHzDyZozK+liNTLGUq2ovmzPzczuqXdNzndMWdXvj7AxU5G3L7IIizDgt+FGAfBNLJnkrmcGK16
h1jCq4nS705YZDPbDaE7fNnqpi3z7F4eSzwAgF3DVOx2FQfUrjMy+w64VmyVobIB4SjlemJg32ZC
xOyCKLnZBc2BUPeHi427fN21/2Jw80ZpdWQP2So4xvJ7ugUE7391L8yUa2G8z9o6DsuGBMBM/AKW
2B7p503ozt/jOvnsdHFiL4yUYiorlxGx+g64KDtQaTbUFQhZNr5/8EHSsASkZRz7P8eQCYnJsONO
Tf93AJvxyzl6X8UFClOigfzQPdVkfkblXtBHcWkDgisJNn0/EVvDYTLmiD6d9vRH1rOjqLky6lpd
77BHzp802tEb6B0NAw+6sViQ3vAAwIkXtTv4A//xnNcS94qm6/HUYMCDuJiBjuoIOwVHPICSalmU
4HEZrRJffAElnCeutsKdtjl54/n85cB5H0dSSsdDuP71mpQ9uVdl3StmcMYRvvq66Y5TztImJU+H
ArVQ5WIJJEo0LszYaNOFEe7h85n78HnLo8fmcrSMc9ydhx+VrNHuJ1Q2j/7VakORS9/PQgf/73i2
+nE7KTpjixc/zZQ8djLd2ZvLWDCzqcZp3/G6sxGBPJPXPDRYezvvAbWU8i7Zaa17D14kTBMevHwe
a/bQCRW+lUuT7Wot0J7qiApOjWyqO0SED1gEefxKmmHfgfP1SKWfxA8KKSC7bl+d2zfqVI0sEZR1
hw82AUFoTcR7Udn5l0nOq4qOHNFwzK9MGjFIOvwCTxsC5550upRwUzPSUX3EaSHSZl4BWeyl5oDB
XWhMts8Ea3HhIhVfn0O3wNo2Z7Rw1H8W2VKhzHOK5/u5BFlG19DYXl+wYpvzMmsyaIfmq6IVtzID
mu76ikGVp1cEbIjOZOCij3Prn074r24ALSzSJ4T9XG/uNtnddP8wqNcuRT6Nz4ORNKao4kQ4RbdW
t36XvKWzgulHbgg4eDLE0S6wNrEe0/ePaU7VFR8n45LY2gC8IM6WDrapQ1E5QfkiaI+2dBpEXR68
zY6jhdJM5RIvPCwfVd7YNswk9E/jURNd/wySoNygxxCEaXvYgsXQF9pgktRPcPDZvmr5CWbxJkcY
c7wbecyVM+hvigw6e/mksXacqXZi6KcoPqd6yzyQ00gzKXPiwKBRHpW4roY549qn9nvA8RaoD6TH
l50MR2YEkPuc/kTmVWAj+ZFYY0QzBjluY109lDDd3vuJ9H8xZ0iNmdR7WyblSW93CMHDFedGqedS
Ugcfg2M2q9msMzG7XlauseIZPpmUagC3Ju/yMT/c9Fjb7L0kQT84ADhSH3/CjW/wXrEf3nHe0tTV
VtxsbMNe9jG3Kvr6Bf3OHfSHRQCpfglJkUkQGr/xSCUe4aO2ljAq9m4FNIO1tlRXVx/Z4GsZg29X
E4PRoXrP76DHJHT54g17Y6Oz828z0rHCZd98QkGlvEdWrkHux0OERgEke8k5btMRVxrU8TIN92vl
p+hHdCD42EEjGO0KI7IuzyfqW1Ld3Jsb9dOOMe/MAxprbj2L2CvbEJahasc8H3l1Uh54Avxlh+bk
4zV3nt2a3XYkjWMzbNDGcVAAsvymBJWxoIS8lplK//sVsmH5XAmxlPMaTrYetyzG9LjRugnx8E7r
u8KaPrhFu2fOQ83ivTLjYb7w91TNR4+kjFHFRJ1sQWHa9uQCtBfkInCRI/D18qg1ErgJGegSBaB+
vT56BwVR7THQhKc1AUD2TOLBcabSZgiJr6Sl/vLxmM0lddDhvJhpaBjObfZBGkxv6zec8cE1wgvs
FVFgraqPqSJmZXsT3fF5QQRPRSxHLRcC3jHSRoyO7CXUUQQYBB5Tupptwy3OyZffeMBqd5ojXroK
4EsS0csmqee2nn1HCsHm6jeDJ92lrdIXiidwP0CQaldL7owsTc8WJtB+IY2PGUmPFYMf4tPmOGdl
tTp+VCAqxwnBkGRnUh3JYfuP3BeJjn6mLzWRur7PdlNjfkO82TqaH2Fn8yAZZJiNCwyx5PjFDuux
IxZdhmJyCwhpktj1Uhd38nj+ATOuaXT0NTp0uhiEOfVmeY9WZPF/41vEqGkE9o42QMvQy7voIdcH
KK8QFGZ+QG4+TLltC6laBCjR+xp53rIGWlkFEJ0bUP6NHhGnYALXqBbqmyszfjmkFTvSAeWIU1jJ
L58Jk2QRxC9jaz2XM/hQUXrUQ6w68Qk6uTwvEC2ykLXRkehnSWZa80xOP+PMfQ5OWoSwdMmltQsq
ir77L63LRrXZ9bDeiXnPKDu15mI0Bx7O3g0jxkkXwnoOuUDlktb7W0dotSjri/bZ2DWTcNATwqk7
xbZrmmo0FbC51kkGQ89atd3mtzUbF7yJzzwUpiBVnSaFojMVaGAK/7Tw7r6RmZ7puG080jvPYd+n
O4LIaLANWUJUSsGr74Y3JCkxAZFwCLpuhN1mZRMaY1k6UAB84xxLKjGjRpUrGOiKo5bTvYb72xum
5DJF0PtdxWk9czecNOJVWM7OoNLg5EiX2j18J+11imoGTqA6c4Wog/eTqxe7EELRhvXjve0qGGH7
kTJ4y5PAooCsMssQxSzmquAWkoVfGj6utnNfCfZbb7xsQUUAUcoKV1mnteuwQ2/kr1AzJErqlph7
UH4I8IeyEOr2RkAJc9M+YzpVwNMb4yz/mmhHzNZEpGxZjiaVt0iMcbCwOjxJgm6cgjyj8RyLRuSr
OHw+d0vmdCtk3oJF0ui5hCokOt5IVzCJzlVCPP7f6ebu1sylZz0LctW/oXgXiAS/oYYXJlcLi7XV
2W5VCcn0fAIIJSNxp+ax40Pqkyes9JPzDW4iQqy3DFAYZ28+n9OcCdHy7UYOE9e+aXkeJgCGvvQ3
BHxMWdvjwkZFGHGBKbIMOpcYo2K7PaeAMyM30yNary20/dzlVf9RyDZbysQEcTKKFJDmSSFoWLYb
iXr0cd4ybq0AbsTaYkTe/kLKP/N/5hyZIPrbeNV6gDU10CWkZmZBN+U+pcc9u+8P2azLhndm5dr7
Fly8xKWIlksMqMr88DbqtTk96lGxS5g9aR+2Ivw522sd5/IZJFZdwl8KPhk/uwOknvVyw3pu765X
vHsMVQsPl9bGyW2yVk641cp429JzLS/zluNsqvoWaKyYMMr/KZII+d8UuRaj54GsulitdQT60n4v
9RTfz24XsEbjQQ9aprKl6T/vWCchaQyO5DK3CLAxNqnkhz8jGNnoQ6jKP4cIXtQ3yHKKzV/eiujs
hdfzkc5MWUplKbeBO3NIDY4PYvdHuZEa6nuk7iAaPHTgzVRokjFRi548yPWtnDPurmr4VEWPDp+2
U3qxYvOnlx/ZJ3cmpntDsTx1CF7XDgbjgwLe+4p42RNF789q8iQh1hAI5lbcUrToEdpkMaMHSgcb
mR/bxCE3WHtHrrzP+CDg28xNoOhBqape0mIyxPYw9Y8+5QeJ2hsRHgtceKjInH3aLha58Km5pwLB
QHX13k3ZSj5rztyf/lJWDU9eZE6Bp+wkRKlKaYhxPKK3dJqdHFrYp55SYjx0YrkkUmKqmOZuWOjo
5qNp1N085z4iTgMj5HUgKcmgqy9ABUCCOCaKX8PwZYVxskjh+onlXtwINeAu53bDOg4VQct4JUsa
M0CwIIuUZsLgTqtY9Cut02pmOOB23GG9g4Xt9xnHtI3GoWCymmzs3WRPhyb69+WeP5g11w6w3IuZ
BIo55FG9+263tn69iSqXL9pCM+rqpy8+RELRA5rzvVZD4t7rhx7uzUz+sB41r6Y2RJ1Wx/vKQSnZ
3di3zkrPbAf4IUz7knao4Aij1O8Ix4bIEUTrpMw2sqFTPouyP75N39CDuv5+j37uF/rlok8XPHdq
kuNwmgjmN1xwvez/E+B5KuBLIpoZXcVM+KW0xbIx47/sRMKYtLVw+T4Q5L7SfEouOlXni/2omaZo
wbvYHOH119G/Bl/+/0SCulR4wP1TzfBifcB3HSrCYVSSXpZu37ZyFLdRXeJLN0O6i8cmgHxQjNox
EeV8blv6uAma7oAvdEvRhr7v50c5HdSJBY2nX5WRQBiAWFBn6P3lL+5dOFBOM+pnqqduf7ZkmBqr
jlgxLWv5UVWjpGIR3BhAWRGTw1r0rXY64h6KO0MyNO9WS1Z+8xukFL02p8HYXLEGTND53xmr2c8W
WhDfKPz2/d3i8qINsi8lNu1bez6TwI3sv9hQ5XCBzgVlg/EhHSp/K7v8sMOZ37nKU7PMf7dl7mUb
dxrAh6mMZPszX3WGjiWQwNDVwjkWAQKpgeZ6hvK/RfgOMWGJE/lRCz//5/xhxwm7IlU3FOyxJpZA
FMPnsg+PuZRZunYpwjLegpCFcFWyL6bmsVAUvsKWiWue1Vrweby1hb5N+CPgW0KVUZrIWJiXqbMA
PSfIVPHsFfxon6zalkWK3oE+kkmEzrPvfILv4PT9tbrXr2RM0VtBT9jY+zq0doeccK5r0jRa2Rk+
BUW8dRPyZoNjo2iuJ/3GmUh1ROqLpbAX8WH1SIw0ubOoFo64wwv1fxQlcGeWI1tALH8iPL2X3q30
I/O+Dq8bnbd+DswDupONau5LUOd11Cso8LuExOHXtgH3s+yIALmVRvZ/6KzQH8k1b1gxjCCYrQHF
DbUfB3RwVSmEF0/ltpl+ZVdZJHn5GX+7icVbFaaNrZ5pWCeHyBtt8JTAMmEsiviqjjOUqHwkfVIJ
FbrNQWLRA4NzFidgJk3BHQAbHOFiB6Tb0Jxbtlca1aHsVcID6bcgkujldqnxiCzJVJLBdMdaRir7
if7BD5EZ+Tmlb2OXKnVkrTyMuudtAKnpuZzgVXrFdC99wiVMFXhNnPmBbdqecduKr6Y1e2iLgxAS
aJKddjnfwds6r3lbagG2qwxj24mKO5CYS7R9Y3Vd6mnxivURdJm/ofHk+62IrMNhC0Wg3z77gZjm
/1OoBugzd3Z0EzGxXhzLPho9It+U7+bx4ItqfKzaEFomNGAzXTwjDy2DSinjKq9TE5SeFqyQU7JV
zCSSo4CxmWtCtZC4+r3Xcr4pEOxA/ARgePaF+vKefe9nOc8Dg1FTSM8EUEU8F4gdJ9gKksQd+9Sf
mt27lsis9/pidJdPRpqsKU0kIIeisGM8WedGUcnlyih2FSLim92GsDFH8HRV/KR4KjYFtlGvvRGi
onZSuOCKdHY8Z4/3Ft6HLH/nr/NCHoZ5SdjKaUnQZ1Ve+phL0zwGHsclDaesMm8evDJS2kXkLPrE
mLC8uRQfWANmoCnVzTcm8Ek1ED9CUgsYHATPmHoZdkPKKzrXmSDYkBuEywQ+r0Q/W60heBHS9BBF
l0NUO6YVjIstQC+lWWaSs2aU3kHGzhbNo2Zg0vgbuIlKgZmJvXdEd78nLiGixBHGTs8PvtIbXAcp
LivSvUZ0jYsrLc23H079D5P7z6jxQv/LCRoezLa+lYUL+Px7/PSSIpRVrVim5cgq1I8nmAQh84zQ
paCQr5RNfvS75IuLPDm6eovsZOF4eQnXdylBpvjYW/P2K0fQGr6oOxb9JazcWsmtNIJHi6XMrZ5Y
G0zvge/rHZQO+eVaPJ1vdm2lXBseF2CfgRUBB1WPezfWcw/A865ioDE+0wEonrnpf0KkDrMWYdjQ
R5uZeP3IV6xGZP7E7HSXr45SRXb9q2n1Ag4qJJQJw8bNY+zVJct1wF5qRgbu5mrAIoGSt+VAspwG
gvKwjsLHP6Ou3VDfnFoE7YOFG/BlrGHjbuQcIjyMtJvVcxNqkBqrYxABfKoDjxUNnd+OdlKEgvRe
QPcdruyZfwwzK9ft2A/xIIQNsg56Gqto/8Gghaqr9eI9h695hI6UF+bab3qY8jlbINIEaHeixPNb
We9TCSLLA3X45if7JY2Lb3oNPjFSSXbPH7cxgQFY0dEa4IlEVDD0I/DAcbuRomR6GUs81D4LgZqG
DcuFiRheTfQi3zGTUN8qDWAa53sUoZHosPruz6oYCR03AYVheMheXSA7y1VRt94d8xlVrqFHafAh
LeHjto8H9h+bxv6HBAZc1h8y6e/hYUBBbNrhkzOki7xeMyOnpwqPUEaxAgE08mfczfdfXNnZG78q
kqB79s9XSSfMsW5IZmL2rNnLBsLWk8++sezznYYpMy07Se5bMI/MJleYKZYxrelPnTbDg8dQ2GZx
Mxkg8qybJkJg+iZYfv1Gxhjh5e6Zs0CnUbzYOxBeGwzkIenIGWR2l5FbzPQgyV1dwn83Chjt1WiK
llZUQgKyT67yIkyoHKzj8kaKjg/80yCBjPxyU9xFMWhVWURb3Sro8x0Kcnv+yY4Z68WKODUEuQxl
ttk6NbSMDWBoaXnneYkSfhud8KJ5uiFCSwnNdIsqLZN84SrNHw1CimsbhFHQDSdcazg3m1rXuSFo
nusNljceVH9OCyv0RIXhhXakOvTiA+OAHm6kWq6G17yjnLL9fHmtDUWelTkgkwQxTIoZ6WKdVL5+
+Gxi6+XHiuJqAw5+FqMzlagBr34T6bd9Z7WzFcUQ12ZevDqyLRjv+b2IvuW5BCmSIH/jBb8S6MBu
NkLgR8TLVYo6LgUCVRaOi9/49ZA76jhEQfZeq5mGsEoDP75wGD6TuvRyHhUDT+dN9OrJrZsjMvaH
X5IQ8d4hKhCse8Z5y+sKvKIld8i0oF92niwE9KZdgztV6+Hsxh5SvISOuv+lDrpEiiIhB0RPm3uz
GjunQv4GL3YCaTPQ24EOFgAm2WJwm5otgK26S439dh6uvhstTqh55HtoI+NjFIT8dGqwicOiqnbt
j50bl3WOlym0DeARlF0t4tcOPeKFOMa6bMTSt0ZvSMHqtJKR/Ztucrc+p7F+az9PBMIn+B3avBaR
zm1jh8qzVMkUt4LWM4yFqae0BVR/GjWwkApj2KcwMBhwCCNZRNpZfPrtbrjzEHdGTMv9hpgY1c5p
Sp5KtE7b9yVWeYqFMpshWeV4KPfCxm2tpTVV72Qc28F5dyf4OO/Ue1SjPP9IySRRTGClZur5RJij
332FneFaAq+H67bVN0wfOxrdHwRDcTjHSfBWsuTG1zGFonuAMpJjif28VTAvcz95vfE99kbE8CT5
Zcyuj1W5/+H9wtfT650hpcZaQkJ8O9p6DSYzC31Izyo+pUAt+mbapaSIdEs+TabYfj0k6wEj65jr
c590JkRo0pOz8ZBzm6ZnDQnE14/jZXCTjylvyHSQHRH5TfWFXcFYIXXxV+c5eCzbDy/EjRf2azbD
xLEdEdMwfZ9Kbwrzvid/DcfRBXO6y2/MeRL+nIUHrqasXyRl1+iJIPVwrI2fETLy7WyLpeQfI6nK
Mg/Hq7MCVN2NxHgpzpRXJcbUrV6Y+qPHyClCyn28yWBDMmWi7cbO/NWGLLr9n55X3gR//2rsZ+ml
GmpWmNLzz8KXCe0fZdlZHNMnUyfiknS7kdY97zanGUpJR0/o00ekaOQHyCeaPwE7G9JvJCFdNwMX
87n71YorrUXvwE/RupMfL/cZgd1xS/kLuwu3zpthpV4DGI0mAFPi/Qc4bDGh/znC09HPv6SvWM71
hdpNZJz2tpmWxVJCKs90IN9OMtuijOWVJ3/mO1X40bHqNPuR3DhpF2im39EYXbHge84k0eKsg32q
0QU+2/8ubSnWH1iA0ojS4yiTqKjRkoW/m/ZyoJhGzpdojr2khzH08bII6+RBAY9hvTVNWdUf4Ke5
g9CIhCFnor59GQkPJsPsvFsyGDZ1PF5G7khAKmPGxwuI7qFQMTV30yDYz/UmdsiFFyjNbjU5hb9q
h/6rLvU/Jejz4fMzE/ksr7PFndxMekuHl6dMg63UA2kDwZvmSyANFxsMsy37/l8U20RU3iI8mEaR
dM8ECpkQBOWYO0+RnwFUssz48gV/a6WW7ufJkztaVsGOnzPwye0LLqUhopYJozgGUSlB36MQCUtW
TLw7oWni14unIbKw3bYwSnJBJ0ApZLzQwEAVjF8srpCD8wsovorCYs77z9yQWtixCK9972lLec9U
QMyGmvX/YqR6SflPL1v8WLGtdO5egiqUWwdiA/zSdh6U9CWG5OruJ222WlpiPavNxOudbSXRP0qI
QWKY6K9y8HV4ly6WqnWodce3hH5p6ZiEKXW3/KrRk+SFhr3z2R/Vb3mzQUieNHCp7UQMzwJyy+wl
PjtGm+mQEhpxzr5V++U6q7dZROvD2ENTna41APNDqwcFN+++iPw0hkuig3FJFsQzGWgi2AZAUdXp
Xxyh//yhswtLRFiTgojleMtKZeunG3D5J+bWp83puhE4VV31De4pgJ9aV2/SqU5GD3Ppetrah6Ln
pMJRrJvN6Qy6b7CvurSj7tsCJ17XgsqEU5peMOT+tYcQxGaOXbTLGqLxu11vA5BKNk4EqrqSuc+9
VjbyFxVo/oqU2PrswfvQYJanPdNiJLRn2Smvy9wCGgi0YGuQ/0bIgVkgfGXM0xain0n1p00jffsJ
GsreG90R5X+J3wyLxQc7vFPd3Lx9TW8Xf7Z/UkXFtDLf/xqtciOpjHhS2bwSP7KGWW4juXSl70qq
qoLeIGJjW2TMHj9z+01FkCX6aEWdhw+DhfnviKWk41MCQGtkwqIRAbu1hZgJltTKFgKw76FlCqh6
PMrEmfVfGVViReEX1/qqW5Wh2GoKhyB9TkuTPL+vwzCveFZv+BsGqdOvutmjVyLicVg8ffNhR5LG
E80iwLj5MEZux0QlO0hitqlkONpWSDf+xHxFvESGJwOjDKfBBlq5QTCgRQPWo2Yc1VIJlzhRTsj6
BVmDaImyhDNOqS7WsxWw2XwrjFmYd4A/75gHhe7o7Cq80NZebx6OQ2WNKd6DaqAO84F2EtGXLJgh
Sv9XfEVJeLdLgJn8E9hRAbTuuAWgAuPVlVJAOE+1wr63cqXatrOo5PoJBbSL+j+6rnkHSoJjh2qI
9zaSQDgGa5l5Sf4nX9jggIhHjticsPXjGNfXHm5VJ/+BljbN/HkE2f8nEWePwLr9hMDgH2n3xz4n
5XUYXkM7CkQeNIL1DrxUL9MYvU9h/oO62J/xM2pmKEvI9hIjoP6kNl+yE7CwBNfWj3BeH7eNjZYX
ZVhdmEykXsocnlrh+c0zimlv/w8NVDkeajg/vBhigMY8zbZW36nOI1E+v1z4w4h+6p7ZD4Uw+2Dp
+iz5njLivnrwIncCPeQQ4eUNrzzyvpGpRk83Wm8fgvUFT3gPWL+sfZIncV0Yav9z/ZfCAuB57KI7
34q7W3kKA+sjB3Lq+OqOA7iaK+zn/2f6Brr5cpokf35kUhzXZjlaFYNFtdumMWASOIdU5cplt0If
my8FvZX3oN8O+BxZdg9VrTS6M82/Ijp9lRBZZTyWig/oZHW2xYjTGWRqltqsUdbMUOP0N8sur+Zm
xsRDYZS0qRHSoQ9hUsgjWM5lvEU8doPpGByuojUuzlx8JtyaLQWp1Osffx/bK7/BihKTAzPYaxGw
aAU5wnq6b2glf2bBd5gokLLI18LbrRf0pRIovikg2ZU08DP6tJsMVr7jZMCYvUXea3qLf9V0j63U
2EksCLyQn2uz14fef484za29K7/kPR7g0xErZh3oZqlOU1hc8dKXTFJC4bZeiEYhgkIioeIdjsLd
KUJbdOH9hZRLm/AMrEy8wyhUI/e1xvku2T+M6+fB7+W/72EHEIbPloFmtQWj5hjgyRiyBcw5F4Lf
ief2oFjwGuLBS/OTpq8GOaGYTGrX38BaW9D5veQMFvx/R3OTuP4zg2QKWnUubTVRj2zjaDCRQf5c
FVzn/tDHgDKFSLx2M2eOlOZljI8xykc1cRUi4OgZ0wV/Fe4aVYbusVNO9DQabDQxGFfcJbF1Z5e5
UGZkpl+HklxdlSs5nquZebqWKvydZNXvr3hwmmKouTKblGTjLMuaSNi5/Ad5VVXJtiNixqU/3bW4
AkaEuKrWHDyQtSuMkRBjQln7GMbzLI0vgvFmL3qI7nXizJxu8c9nfPjj53MrnBQeyxaso8zh8/1Y
IwaXuiyB3M8jyMxioM2NRN0p75jLWFreVFXXdNXM4AlMZoqil/EIKIY4AL8XwwH3AzE0EyD+v5+H
C4lm+H0Dy+vwxcbOJVPEmiS6FOIx4pFkxlyQHWoIuYsVPmzLfdlUUp4rpXjrqqt8SoDlQHIbATkI
JxoZB0XvBIIIXtnkci1QlK7I9daGSAs1DOhQ6oYKcFiooipo9gtoka72vhGqqOJ/32AzL9853xwJ
+0I8/owQD89R1OrKMyqIYL1dtkyjPz9rRVYU5lwSaUGlo95fYk+V0zeF8+PAscoQQlm0kt4zESlH
/skoK8VyspsclENvPWfdnsmMH9kJ6mHI5zNCahARFwNYohPLvP9Lwc656XdJ1C174NAnbbB7yAge
BB2KRywyQyQyjzmdWPQFYcresqbthx0H6cxD/oqm6USfgvfWU3TIFxUHGyz/AlwY8YOCngJayGy0
4x7OSX/dVt9FZgH17jsXSEbv2i5eWJmEnjBplk1+wIJM0Dnk8XvwJiavUDv1W4hLLNg+wgmSPFy6
FyyVcjjbU22WMWU1+J11duzc9u/pBG+CMMjs9UGqRt+GK8PAyxa8/M9BCB5wiAhWxZW4ZEep43t2
gNQz6Ct8agdQst14J7/Zni4FjOZAovmN8rYnwoqjgM3kLDhix1VhssuRx8EKTcuQ6e+kSHyYsyXF
RYTgroncadOJKHPYCOqmKaL966OrDNOR9gseuKdkshWx0VTnZHo6P96A96S2a2HhHud6PmqSAs++
t3K0KxBCHTqCS+S+91PzEvltwLNIPQl6qakXK2njC8bW13nUPMTVAPGopMMNanqHciMuaoiVCfzq
hYCYueA4aiYj08Y4SBgieRgN51PobNWVUnsnaz1cu9I2LXKWz/kfUwZluGfS1m+RdrwwFvh2JiQ7
i6D/0KZQ52/Xassv2YDyI+/dz0tdewmnym6s2uZeuD4uP+VWgbx/zKTpkdXIXeqRBzGkrXLtORTO
w5Q2wuFdiyUDS8vvIjGYheNfnKPIYOk1jFOOdIAz+/HLTu/1wv0VRa2Fe9b2tlPnE0AyYYBUqngm
yWYtdfcasC5YzLb1jurti20ApakobKPRzjVQe4nxOFU98D+a304L9NqmWunhN6utSu/ULdSRSirI
2eUn/8W9el1w1yS4sHQue5awAMO94/8z2+bn/ELcNzECUAVvvzjEPksHrEhUpVBkSuXeG+h4zUO2
vY43XNgqx9RxKjU0Kefwkg71G6Pxb8V4hZjAk6o8iamIqmHP3vNT3KMWw3X0fMJthL3/ABpAIT3o
Q5Tg7OnQ3Lt4a75VT1OI6EobtJLlw+AicJCZaC8iJ1L3wb8OjY25fBDaNJFWtC7qazkUx8PZgQZt
tzO40ljoPZVMfTidsuCz0t4tKjFUT7sCq2GinSTBb6qJ/ubUAEZtOaINduccPlU76w1xk8+VUReL
yy7jSB/TJ2HSQQWhAJLA1dbUKA6aWZ9OOws8sO+r8fTQYoo+DbgMRO8aitP2/VKI4MCu1mtiyOU0
dRkxp2scwh9DllIm1F248XJR2xoVdHHpqm029R4xs0+735gyano3NqZzJFb36cDoMsNWQUhOG8CC
dxgT3vgmPQqkgamRftdeSvmk+6tYonSXcI1jWy2DgQYGchRRXpi7TlUfIMXVMA6HA/1RQNi22vXb
mWi3ajQQM/Kot+b/l4qUjE3tCEqKCu1ZXcElrfzyVjjAnIiTXNsZrMX8VdlX62XtXdKYoqh5nX4N
X+qAroeMif8YCHg9EkaXZKp9QQAvqFrsocnX+NAob12OJZKHOjy9S0x7GOktlifquTFO5DRuqrAp
LvRD0vmiO/WRI/q9Q+rQ13s6+Uq+lJEOGDQXdjfyTxIzHRoYMJBX314MrUajKz8g9P9k/pHYL/G8
+Jx6ghDumMrMLu7N5s1OZu02T/h9HTWBgrLR724Oi+riM1szM/hGUV4UZ4Kvgfd14ZB/qJJBfKG5
mx2bKWsoHJ0JNKeH4lpOKcwj0e3+LAtK4uldymisdBcYxeGTE05AON8uY8FxK4ckDQJ0K/0lXmr1
yZxIzPloQ9r0ZcMgY59os1TJZxsAf3g2UFq+9ejD5Qm712M48UclhaC10cZ4JzXvfcC/qcXGb39o
3Pog/EW9op4N+aAjREQWsv2olu7AuZ/nrAWIi5ssdWVzfxCMxAvLt64I5m3MgCFzbyIso9Om0Ngu
SgKf7H419a/Qhd30Pil7aGed/G3giJXIP/tikNWsxGoqEBO8r0K+5jVGWyWMhUaemQpAtgYTZQGq
RtZfflJP6FWcotZZ+FffIaPk3rrlD0GgaC1MjRD09XDV23JfmypghwtaxnkzbfS3tiYFhukMRkBK
TF7/YYsTlzlAFXDhmAXUBUREXD7kHZLzlBGFKYC2SRZjdGh4TrH/IgsaCPjlCwWas5tuWmGoGpTs
Qw1Z5rut6HVqOwdpNSvAVei8JWvc3olYThuKvMUHo8f4shHCQzrsNM0OCa1RGvraHfi6aRcM4MDf
7BXvARb2KCPzpNCoyXmH2Hr92c94swEr+mSoET63vHCCN1ojrkI1p+nopGPAJW6udPsE1VeNG9Av
kYoKTSK7X6XVmX0UHww0lgTaPAnpEy1o8WMcdNA4GNuUR8MQCqtMdYaaZapv5jHehZW+Kz8RjvNu
cPIdZCp1CgfwCJUYcEvm023dDO+/glkKO6B8TeLGjxXvm0gSb5de7ys/sxc8nNoXjXcLZJP5SFS5
Nw3+yXiewotNdRjYq+oF2Qey5fTmBiB7Co39udHYmBixJ1mpeI+6fqLt6STcvNWTj8sw/s5AjjN2
bN5Dsyy1UFEx4r/zkMZH4VtTbzgi4aPBkt/MdJEop4UkygTTYOUL+5CUrBIubeVf8TU8E6WkcrjX
MJ7ZHLR8kU4VU1tsiCDRtjx6EpwySKOKBd97BNjW8kScvoDC5wMjwR9bM8ATVDwyMGHFkw2szXR6
BC4fs1iIKjp7WmSJV5nn74d7j7JU2Fes5iy1pJjOr4y1biF9SkZpI6VtdojOJuqtWVuz/oEOaTcN
xMiRXPLvDRE6H/yi52+rxnX6TVCMVxosGeuZnCTohPM+Ts+2SBKeqfuNas2yz7TXLhSjnZr6ez/l
x7SKEoNJVLrKREAd7CAXwg/It2p7H53c2+w5bkVFz6akpP9Xup6GxmoXlrZ5upCjngZZrAX6rZ/U
slzGcaX//WylQm9CBwf1fAcA8EFOcdqPt2fv2K6q+GbwFT5Zvc6D+N+jhDsmFr/PaZxGUBmlwM5d
z0bKJlABX7U1sgwYStRc4xCTXa5UPofCcKZo5RWGBpkVFEzfB0dOLqPc23iphjh653ncCLmi+C4f
hF+zcN1w0G0P49txyxzdViUVkaKu12Ngdpckvi4qb7CbgAm11JN5wTgt9+YI6VK9mWnEkhrgNioN
kOFdtb+bSUmlyHuV0lRKyGy40kR9tAA7UasuoNvUzOWmWQwNa9LbYpVAN+CJIlGTGCDRUbgdlkKQ
MUbz4rgsQfRgi6KDSYfdlP4xHbxAx9BarW1HvIzWHTLh/WLNjEDYQbOIIAdvoc5s7su3Zh6cPSEc
qREX/D1E0tYio7tNMJl0wpLDP3EM1ow/SK8S0Yk7dTSDUbCu5wAAntL/LnVbIjaPEzUIFrXiRi+z
lW9h3QvHRvHoVQjdbZhgH7LtXOricqRLbmNJ/Jupr0B3FnXked0NGYyBfJZSfObXSRo8J2XSV5Jz
FziYLUBRVN50GTGe5PnNSGRo3HNhd+guE/QvPl2d8s09bGNHTVAL8UCpugNE2obPU+NawrLvzP1v
Ybg6/9wrlGwzlEL5u7lT3OdR4N3TzOYT1ZxYhwhR8ohy6xVjqmXbwyN9fLOb95tsUhEICNyWS8wN
2W52fMZz6rIuYUmRZ6Tia6W0OewqQjRC+nD9udEtPT8BMj9kDGKsoxo42Ztpm0mg+w/pYGMQKIID
Gj7YhxaWUKwNuXKZ4fMRBIt1ZpJzFGEXbCp6UeJZPb81f6B04qpeepdBWp83mxk5A+e7/ben9XRX
CQ545X98RFRx8byp5orQZY1V8LKIbpBQ6owM1Tf/8QXICCj2QUU0TWFiEiSNJ726LQUuqeBduQoW
hSrH7knM3qXV647iPSGWzrD6cRPDbgK+RUYcPmTw7IyLpi8vS5mDqr+CkSfLeEBf68doBVZkal1K
DyHq/CnEwqIliDc+0AdF5j0SuQUk1uWLxJkoYpzvF2W0nvbH2JdyMpPt04aC1PfIU3IysMq2GRJS
OZoHyaszOAeKCgtKmNqnBZeuY42Rd8bQA7aU2UkuDzSvZfurhQLdCFCjX23U3iyxg4PehrLgMhEO
Xh1i7pP+xeuwGuQgN0mrr5aie1KnhC+O84AjYvBhEYq7aAw2O/JQaa3DSwOj0mTb4cnsx4iK3YZi
FWgrcnxAWvmy2FtaLuxsnOIhU2/v8X4+NChw0A1rovsKje1fYWZFr3R2yjyKz2P73BjoaywUX2cP
75RGovuWBAOru0+yUnXCE/1TpafHd/qJOmnp4JSvmEKRsydUvx2/rO3vc96SJf/QvBtAn91d/Cu/
jkRs7qSgjabBIajNNyuJzFNyNo1XpPcIc4zbXF0hv6q2GExxt11bla/UlNAzIckAWLdERPCTjj1s
MEeCK5V/KmkZHqGjYSA/kHcuCREH7g0GVOiRvkGFLEvQHdaS+qG51OFSNLQDipbx73S+zEhYc5PN
zMDJX1deW82WIoElPxKjD020tTRs/xWWwFUnFG19gzK9tycmtvTgZK7KJfAFUGFv4UynEM+I5F0i
Kv7zANnhFI4o1Z7/RnqST9oXFqx8ly7KbH0siPKJf8343XOo+TMYoZXcVxpnY5prZGEZstK2ty8H
vdXwDAMQXT4r/cCauY+nbDo0IaLcdL7gQlIWnAwYlsFn+SrbuhgsfuB4m/QFvwbVlCBZyUieLedK
H8x05Iw35mdZXnQNbpEHuuBYCg0JFm4vQ5OJgp/HyvLFHd83W3mGvWnTIXV+R7d9VRis1dpRXAd5
KP8ve7T0Ik5P2V+dNxCgQOP23fe4jeyqqUUi8aedQCkPXVEenSGws5XuhcktHtAQndkywnqZkZHK
pepf6CKC55jBRuNxtUf46daH48dC+oCw2uXJU7v0K15GztwbEK7/Bwqup+ZuPx83LOqaUMztEZ/N
BAiugT8vsHCgcIvjiP/ZbfjdgSFWUG9eCW4RxUIt/3BIwbpRteBEX540eJecxv4YijnLiCTQi31i
LDNZDVowL2KTUTBid7zkUasCqNdGObutM1C5n7TPlGV4d+9edqP1wzqVy9iVhrz7M0Z7ZGsJOdpf
I3+kEIG3qqgv9iw/WX53KV7fL9oFsU0EF6XD2SsAoS3OFwdna/jV9QcLy6HGaHX/YMGwLXzF/MgV
Hy/MsKqev2lZ8dbnyFP9pySxj47YEIqm1WbF43DzKkcXs3kG8ANx5D71Mdj2F2a8JA2EPRa+5X74
6TMB82ti3nz6TZyt1VdhJRaTQKC1oponOxR5jP2deijPBI3bz6K2N8hlAu0a7JeU65ULfNiE99em
ZLYNlgU/s7z4BycQoigmVVN+RV18m/CbTl3/1vU8nDgWxmyYTNOykRZ4NSNzkVjay+baDxfax0Le
SjhJomfWGl4dfDkq4yQpaZCR/AOa5F2oYu9PtYFWatDnFePLCDPeaVqST/xFTYwOuSDr3CT2BGwC
VUVsqm1NFzk6AzcK+UyGmJM+BKQywXzZ1dEP/+2DKQs4ZKi/gncdvW/85I17v7fd3ecPvpRRXg+G
QJx7M5+R7CuYNlrixba5+kGyxbGqqG+ZM0P2ahKXWHrOsCxEoo4MaP8dB5yhQfYiMJtJSKGgepl1
R9r+dM4dKoeyA/cITqGv9TdwdmVC/uG6pap+tg8fEfRfKcusxtexc+l9/Ler9CMZm0rhAEPkDQiP
GcNX1ktjvh/fQG3p+KAnwfdorEr2vJl/ixlFqEOtvtqaobkz3BuxaMTbYm7bRClhcE9XJQ19qE5I
wPIXOXFtTTojIOMNsMWJPk/Ww/GQYlmcKMchvF+sNAhWySNzetl1LtEn1vn7is9Zy4jjrUrYj0Vd
UVhFKfKQcPCgbQCuwpqyhGDazh7yP6cnlQfQXiXJt8KgrExTBMUQNYIc/kt2UVp6d7DVhAwxjajv
CPis37ySGzdEvyJQugktm+wDDhPU015s1YVtDjYBWFtfQ9dlWM9YPjscnR8dh3fZVb+qGWXxYFc9
e6lDXpG0Mf4XhlxwpWRXBjXestp86sIUAaXJJrpcILeWoLuezf/26ELQ+xDvLH4ojj1zMW0TfleS
kTbme4RNj8L5LPmnsJzOxMKadM/9YMu7xOSl55m42G97CoTlVmK4KpedmFDths7hbvwCWRUeE1FQ
f43lSWQdzwmfI+AsaabpHNpoj4EJ5hqxzkncpcJfNtcNXTOuNC7ZnKnJZFVuU20X8Gh4hplDLh8L
SyFEeuqmh+DywxYhnVpjNeNLY6Izl7xHWAL5qMLppe+9xBWmTRxmQJ8Dlo5XvEhQvnCEZgrS71l5
z1LuFir7n9qn6OBTZNT5uLEmGyMDqwwcf2vj2NteZQ4yKLH/jhzqG5xOA+kheN+btW6MD6t3lRzZ
oJhJoPkEZg4QnJx8j189k1AGROOqOMsmViAA5YT+t6thzSON9uAgCBHND08V1wSwjDKLzMVlJ+e9
/5dYoqV6gsh5+7iQ8gLzxJuRXuS5vEZUqLIzoojkIIzN6hNXuImFpQJKaCCBbdnupPSrH4CZkHXX
5Jf/Fc29IvRVyUxZ+Q7xzPZt53noBChYOFHP1eM/IrrAramr/53ri6GuI0blxbbwO2p+dvui7q0r
g7ZyfIuCV2Xlo4ztIiyIWJWEnWLcazUREfDNgiTrhV6P3UvBaCaSwAzksvGjt41BEdkODjKjFre7
KpXYYZkSud/dxkW8FeAyz6AGUqVugGcmqSInxXiPdggl5VmYPpS7JRtxVw6YkLdYCbfhrvYKL57j
m6Dg3ibsKwiisMi4WnsYQOue3WRdXoJ9O0LDORRtZZnSJokiMl6VWWAAsiXf0gKry76/ld2/eK7W
IBl0y6X5dhUXNZLqzKcBYsohHfdfRjLWwpX1OzLiOk4OMgs7OTuermCGkysrKRcdruiDhCn+6Sk3
psG2xkawAa0Ug6g1Bd0h9NbrZVfkxkB4oA2vWO6yyCIZAdejow04tG0JCjyLFhTh77br61e7BnhE
oKfGZa0BmG7oIDWH2EB8T8vm+VIGdfUOgHv3OLcf6CoBuChG1XKclhS8By79SQQC1CbvMUOK+xRU
VNihZFFwmQHmIBS7tSgGNpIMQa6coUISzdQnYb+4EcAke/nFApVeB3+nRKpC48JB8mJdP6jGHiJf
VZ34ShY9SPhHtSW5oVr7w0aT4MD/XRVpteaS4psYg3zaQ+YjE1JDKm1aGtPeMiUFKEu9If9UO429
Dzlzt9KxiMG8Rfn2wH6NDOtHcfP1j0Dd7VaV5xQ7y6UPTDx4OoA3py3ebb+Lw55fUIPXyr1AOvIH
FLmhsGt0iMluYgNk0xO3B8jLN9womDG+b6fVSZ5ClG8XUBBG8nSOlfVkdQ397dml5yaAB1vGhJjO
aIrelgq89OtGRIp1bcfZHCGXBm62gKxuLot6+a9E1ETRhCssSDGfFDv7sv1Ugj87/E/SDjEjjJkr
KN/oS+31lOpOu6zKFyml3n2+3Dxk6Qp5MT/+imjxCXOcmjpQKj4YxLmu0h14bayKSVpyKabEMy2I
+lfwSPt+VD+SAne7RmEpA+G1i+e5LbR8qxeF5pqFh5WeMdGMIOlpGOHoSD7/IgEGT6dhY+iHRuwO
KD+hyM06G0hg5sziQf9vDKuAja5/Z/XtxKA4GE0Y17pYGph5a0aSpytiZxzcniYj2KPzYocLxRZ0
B69DK2s0s881rXFLmx2R7P1uBwfEzzv3faIP+1b2qdxANSRg6h+fGYUA4twtxti+JDUyB1vzlQS1
AzLNmciMxnRVNSRJzpowmRYI5Q3AeA7rQ510ylSyR36in087bGf0QQFTNfU0pC5ZmEKkd0i1Ifre
nFyfYFU1/B6JJtxOoqeplXZSj9G5Wlpqm2DhbHSOT7RZIJ8LGrjBtLiQX0CUUzh7OD+frkqSOqqN
wj5e+TiR9aXBq3WqsspoWgmFvoeyONXVJga6qZITGznFNLGUGjOgaTq3tWzNiair+1Q2vjBA8AAt
aq78Y+yrIGOOu0FPIcc3To5P0EoRc3E4/EllYo85dkj4Djv6Wq6WmgGjCbUTZxd7J3X0Qg0tQ1fA
narbu7cltv/s6Gm6O4iZcrgPX8Kd/9fYuknZyHi/gzoQhBLgr7fCfi6RAh8H+9LQZmhLQT5xauuK
b2rnBAi/Oj3uR8AFaBXKHzyHctGi1r3szqF7RvjNQeLJbXu5q49l50Wy7ZK+TJ4hEXjvD2xlqzti
SieUJumttOgrBvhMg2B+7RTf6WdfdBN0fqP3XO8FbDYiorQ8kzcaApZg5RBzSIw4lz8JXmYbOK72
RpLImqRoNhCMGoIsHzBuixxxhkS0YpGJDMSI4spNAR4Xl4FjThThPeOpxSVX9vWmYwYlfDaeoHpG
ElUtbETeK+EiIF8aMJaaugK3yDeQzGvMqeHO+4uM+qPKaP9R5tmgeKLVoXF+gKlAbGnxYjYPZczT
eEpHaOEuX72tY75byp6EFPiTlSdjIkqZ1+eAWrlDhDvBKSjYC8/sg43SaIpHXDem7pB30yDdRoYr
3PmMkExwqL7m0rHZE6kYW85/4QeSMHPU337Ime/BaUR3E+mssr1y8t6r4So84oEjbBc8wtTetRsd
Yw3I8Ffy1BsXVwz2eprzihfURSynsT66TqsFnhFMrPcBuOIS9RCeCx38HxPOwYZFRa1b4CdgHhHU
us3NWU7bHIR6RxUWMwWp/CgK3CkHL9dLNzUFIZ/7MvHAqlzTNaIgVRsK3e3NyhQn03MjZaEqysem
G85zBuaXemGP3rMzasQz85OCpPsc8ILb/Zl6gmG510a8u0xNp54IGrjsTBF8VMvXtoMbC/CegAlS
dpG2RHUDwaPeIwL4pgyplk34uKbDRR7kT4s7R2NSpuhtZ7giHjTPSZJZRsiuXhs0HeDdzUbLuaQW
Gjav8w8bxvoDb2Gm6nq/8KOWv2wDN1SCgLppHwd5U3chMLUv7blKheJ5HGPHDH8zYQTuju5t6Im8
V0bRdwh2ItTYroqnTzf85bv9PzuNbzwI88bskmi3vcjRMqW7marxDZ3nGP5pbzNEvm8QYLI/sBEa
sk82vNffXBfJ8kVn9nESGuhSycMSoJiRGGXMFlIRbk57+22tbL8mH+mVyRo0HNT7sW/f0czfimqW
mpoZ1F76LnaJ64T58qAheWOdEOT563zYsr8opO1A+r8LQ7BaNVNlUsXnGPAVQTpUFF4tZSX6p8Ef
7q7OpZMUZdQSPrrz/T8macPFqpqNHIavvdpfPLWIO13R51rtG9JMfASyDO55s+7rkAT/8Ay3cApH
LjlPwuw452Q4x8vqYx4Yc3rgAYDX9CUHX+AOgE1e1oFK3IoUpxPGA4NjNVhP3lg4FWAzjIiVzOae
1oe3EzBEyN1ODCyZWa8L4aJ53mK9/luzAw8G4PZMwBOAjb3blG4S2D+EenJiKpr1AJSwlc43h99i
srdSrYDZpxO7c5EMRzougmR7ZtF1lg/31fGsBz4pvY1AscySPPZdnGHxC4boTs5RsH/mqtPj5t8H
Fn35/9F6xIX185E4e/ukKCSzMDabq/2fkygLF/8iGXxsVGkzxtOrlvoUh2r2uutLRcez6MvwONt9
sFNxdwmAJruIOYInGb2ZhNIHOyWqI2IeOJ7zq68SdkFiFjrRc8MHQ5Wvj8TcKotB0Ak4BXfMe944
LdVY0mvz6jBPEYNDBbA2drcOeL+rSSf78cCV1l/ir7R0LR1tDImXtbevemmEIhwxj+wUyymAkUe7
tsYRaxO73pVp975HbOsKDOksdMQs3M1lOSdZJqHDyYdot/vCwrRPV1FVSvffIJdbnoiVZxEnNcN1
yGqAgSyCs963olDngVykgLTsR4tjFAPRwYo1A7n8LRnn4xYekLOSlCguSYLmfvG+XNzgkT/LgQyX
Kk0rydCe80SKZ7+iDs6KySpGu7rQveFAanCT9sXQCm58rbXiWBf8VZpDvazwZq8EsbmDberQo11y
iS7F3iBg4aEywFbVbNkSIG/Gud4bIP/gBaOPaMLqulUtcY7GZtAbeuBUgZQTa7Ppe67XYOoWqOGo
ijHeiEVQd6/fjsX6wbjoTQoF9Js3wAq2gktlQDI0ppUeITuumMihWh9eDWaJs2ZdMMZAEvwI4BJn
dFjLebGqTA2RJFuvReWAz+9zppaMGLaUOg6QgILZbwCbWKE5EMa439PfJuaWzWpf8Mvj2mDYhMKU
1qU+DKBBCsdrTXJ9uSvb3I4595COEMf463aekiWrRN0LdXg6wgB/HIKNnCPbgvkhE1WpMinv/rS/
dYaXOewSilGta9M/qcYUEb4T4Cbe1Cq3NVE/frxxbBd+4N5663JHxWUjdLsp0SFxMztjHVL8BYp3
VQpwytswOgshPAF83oOq2ffqSONl8pVwojBTYfq0iaSQtshl0ltBUasGcsGmUbKslAb1OzCaP3b0
PXEOv6m5yOZ2WxcwpoYUTrWjX7D3Y5FS5i1MYadv8xNy1v3PxUsLgi9x89dzx9QcC+AqXXhJUPqV
1N5lzOUtnh/rvqIL9jiXJt/mo/8PybZUVIxEtZ4JKuw1bcgMyzozmld/H1Yrz+4Qh3xdmIvWdvBH
lXUntr9eLf6n54ZoDadzrB0RuqMXhzxEn72IC05ynFnB6NPXZZwFJq7BeNPoDjYdlueqxlkjIJrz
m6W3Ba8/WAGmsIc3Ky2lvjje9aqbKbeZ5bW8GouL0MMjibEUALbwsO3Yd791LuWMMp+WjPCgBVwo
Y+qg+I7I3HkNWrHxlSNlTmituDQ8S3JWfKQQoS3XSXmna8cu+eOQ7OWuSLlevgMDVH2hMG9oZO01
BRZHfjGpbUpsBQj656QvTTBfCQlV8Qn9MZEcmsGxcZI8Yk1m/K9BY3hWLBnUPfUG36yIpu+AjL9e
cdnwLs0a8HaU/Z6HCqwEDuhk4apPAklh2pvTs5oeG/lL/jNKwXtPP3KF8jCbeCXlfyRKicQt6/x7
SEu7rMRXrCLeyFZhmIVnA0C8F76H2r0hn6gezyDx3BAgWljReGRDqtTmVA9ZMEOMDtEB3n81I/pF
pNxXeFbflwfZZMS/i4O0ALW0+4DfvNwnHihFpqYrbWS2W7p1seuB1ySeB1WQ8cLUFQOKIOwlVTEh
EgkBXCYDXlZlcpef9XVTefxwChpiCGYarCV0XicUN+JbNJk760Li0AvgM85eazrjxRP15vLCJyjP
BF9+j1v/aaZApV07pEFQO5FXsHIXcrYY4cK+oJ8Czxn9sjXJOJAnjVY3yfbCN/mziZKmsBCzNO8P
B/VQPvvcDe+t8rtjHgQGpwXaQNqJdLkr+cj1b3QCxSK7X9clIBbjvQevtO28xvNQG9NXIDN+PBP2
67/Cai3I5b9g+XaRIf4N2fzrWk1CRLTK1LoZrpP4gOwj4YEwP6g56VTGqvK8eUVhklPj5zp9Lyw2
FRIAlaDq6RT0i+93qojyxuynMvY4tGoM1E7wDPCrz6tMr1Hphk0fDjgRq5lLLl8kDdN78qRE0Gf4
Tpdl/D08sO9uzCjUO4ilgKpE8P+yzZz7qErYfl55Wu9+Sg/NiGgUHd6fnV5MlXfCnq2JcKcr0k8n
ZWc5ZZWNPYANXc3N8fOASMLV08i+Eb9PFRxD23G2lN/NRTD0smncyH4/MMCb1X/CT0VobdhEjWZr
ikQQEwqq6FMo34BbajqOeg+fKE5nIaYHE+j1J1IVXE2kaCYwzSEZIFHlmrIP+Ry7N81eLCOKOBTi
l7vN1CnkwykVZ25ztVcuMSEBPoKIfFZHY05g1At2wBm7v37xKdb3BGCEhTi8kAfdoyfTMeWRZVrO
BVGwIg3sFg/Bbf9c7duQRWBaoWKy8cQGiGywHErJwRZXJnq8q/PV240psD3W+UvCQwBOoktnTsc4
jzudcNChSPr1VtSPx0AA3vK7sUxbilkUF8RrSxbVt7+0R1MALfBuUaO73fhBJFyXRIO4rOCdHS9Y
26NaRAkUDgtf3d4ZY5oYrLTyfapHG28V3GNMlP6lx3CA+jiIi/cywZJW8+dzl7hrbJyf4l7az/yF
cDMTf4efveEd2y1SHBbUHVbg3dkOT89rutwqja9Z/d20DDeWaOH0lLMutgnMg40wbMlCbj3G7V1g
1G9vEa7u0P/juHL9DbA5+IisEy5izqED2h4vkJx5tqClX/jQcsD03ahQITlS5yJGObQYjQDB/qrK
lduz/P3utxPb6muUK+pVa1bN7vNQ/j5vnD+r8sEN1Oc4TttQKGjHdTiyVWZd0Ks2hHLbQu7MzG17
RcgG8ysUVtuk3rKcrBGlFXQcyM/Dz97yWOm1NGi3gmv8E6y+riUhFKWOKXyj2nwLPm6Bx4+eThGi
2oxQ+X39qLtaAKF9SRsBCUT8hrJ9mJ0Z7gNG0U1GVlF5aI31cOs9bxG75Qu2puhD/CbqM75Frsa7
tgIJt+9Iv+GmOsI7jm5wfjdZ4HSrTbzXjMFSiu5/5LvDxnhP+PyIdU/JragzE8mGxf1jfOl9tNtq
ct+lhddzayd/p/qVa0eObZqKj26KPO7BBq0n/JR22yYGWn7mAmaxySmjCZ0YIjJQ147LkFpFYIgP
yVNz/G4cRGiFKbmRLg+koUD/hY2sc4aMnEf2EP+fzr/cWrGuZcH6yP1/4NXAks94AqEQseUhyLI9
bjJ0zCwqo1NU7do0IJViFmSgkY3Lr1E2Ildo/DKPXq2B1Y0WLPjVdx9Z8AgnPu/sdGp25cI5V/X3
Nd3M+t/WN8mtuGkzqRgixLvXYoWmczikuwJTpvsmYOgIKZtky5rwWN5CLXvOMhX+3aP/hwWp455s
7HuotNrbOrsgzjCRvySspU2eqJuQjmSuJgCxspOqjHP9N4bw3j770Prah8lWbqXA8GF3nHlwf7OF
TqVMATCFMFu/7ycIOCu/wAW2sQDHtMcSSnPSZ5NN5j+0IDCws8EbWHWYCdhB5X1S53y1dCAYyMzZ
nEFhIDAjXO7BFg96WRBGRUn3Czdx0SW9h4k8lq6XXsCgaLhIrZ8oxE0W89ql2f908Anp1FGfm+rA
Q1EHQWAcuDeX4c4W+KA/70UbUf+gMWdMq6bNHbsj7jRi40q7XzUyPKFM+5Y5sqEm9vAPlGU6Vo0a
GmqJyuCeQmpsuRTgphgG6LES9NUpHJhEIUJBneK6o855zs5yzkYywP0p5P1WZAl8o26cNcnWZe9A
6mg9q1k1j3jXftSyZPSWLbsPSCX+yGHva0cKOVIzz7y2aTVaWMUt28GrMj857tZYlw0Qgexb1gOy
CkvLg6MajrNuUQwupauJ/Znij68b0avMRnpvwqW/CFGbH4bRdCb2gC33kc9HLYt088js0ezkGIt0
g3JxJJmoBO8tp0Pph/1gSYKG4GI9iODpaSm5fey5U5qG1ZCxXb7/WvZjriK1P7KVb6YSzCPyMFot
8R5c7jjcqu8LMUN9JZJYAV8li4h9OtfEjHrhUpJwgg89di2VrxmXNfXG5/b9g/mjsXvaVdP9+m6A
aPnEjZqqsX2SaapBfsiHGouCh0r+jKI7r6dx0urHDG3brBvrriqhNTrLODxmhPYGJE/ILKgI0csE
5mqEkvpkfapKadXfhxFGWhtRzbne3ii17eOhqB1qpwSYCudTQJkVG+mCI/WvZGsl5U/8PLhtM5+K
VDbbQdmBOudKCGyNjmcylLJxMnCKaytwxCwS+yQiWBO8Gwf+Wz5q89cSh8ZXPpzeTr8SGm8USEvG
SwgD20y4eDwxHdmkHMg35B31E8+YikB7L9O4jsZffA2m0Fi2q7fdZnqOcDVBn5OCQwCH/2PPeaq3
8LUoIqc2A1NnOVmU0t4GTjT6DVF5R9EExtwuqbzPKiPJ5fyc5ysBo1/qoid3m+pKxWIHa6Yj3IW8
jY7yzJyqkDgXPaMWP7JB00vXDnNHRl8fEKqNY/ZzjvldU4PZo7EX6yi8MIvDv8w8YFdNqVYLJMtz
i3uKMbcF86kZqJ5drCa2BY/0rf4sTvrKRXQC0DjwWR3qBpVj3sldlYg1jHFIXrqA3tdhbqjwvEzT
1kHiklig4M7tMyfuMngTXwLKyDZXTwN9HQzv8uyx8/EBTHxy++/doWvXz+ECzPLPEUMxfLBkcnQC
bJyUxMtpe1QwM3KuzbAi3KgMLkwKS8rBSBq2DHswLkoaY5PtBOB8nMLpn0Az2CF+PX4RHBffcy4A
HegeSdSHglF5WuYboHqSbxwrdc4k7acRDoj+X2Nl+Qc99PMT3i+HK7fRtF4XkAj8abvFWl0/6WhP
IV871CQuHk3ekqY9Nb+DrZGEAYaULPDS8kHnDU3Ka+HC15OBEgpSj1OJPN9w2wHBzhF3EQtAsQRG
0eAcB2nGaKW/Jsc6dZnUNEeC1Bvt4uhAn/+vvSOoHpVOorlw+en+cEkOll5SF/7OOx4J6I1+cBD8
bT9OvaWt7Lo9rdLNrQBtGElx7Eo4iyzoSgruvfIVSqVfDl4vbnM3k85CD99/JcAPn5zHy/YnN9Qd
AvzRYek26f30Zm7xPGTPy/cHwwV96BEepzZIF8zXzeMFC/gu0o5390RIj31Ezh7nFprUACCC0pe+
Xv/aqVfyGb07Tp9snKUzmR6BzYcGqJtAyfElxyU2HliXt91nz2itPsQpGIctN8o6q1RuccnEeK2/
uRvDDVx0GA6+NF4x30UxBI2D/zJR5dwf/DZu8gRjm9C7U2VoJmNYmmNv7UyBty7SjWgsD77ZKa/8
HDAuGFLz9iHuj+B07mSl0bDBKepgGmgNMX6s/Ta+NCY8/2QwO7P0t4cgzq0HKv41kBggnccqDiHg
1O/GzamSpYR4p1IbzdPwD4ciZDTNli+75xDfZBrRVx/A3LN68I2YPuXEkUi1jE48Jtg6eV3sQF9u
X6Y1S1/DxYj7iwI3U1frhkPzscU/8hzrh1ci+vzPqo1uJemXBSeLqkQOay+LHmjCYegodIHxmBUS
YMPc0Hib4iOER3y9enpfsjOKDfGjt7Z13shhUbjMZhTC553sGP/4vorp/rvzmBSGQAikYSQKObSa
OwiBQN6Kjt/XokCla98N3DxgGQ1NSbdNnmTma82+OSLB9PCho04v3odFHLmrZ8J99hVt1e5lK5z4
7QLMZGVlrW4omNLS5EzCM5so0QTcMiXtFaXUuzjvtK7Or7YRY/oE67kmYEZFc6ZwKaWxiCe3c+iV
rSs/eFGrD/NnUXCRi3P6KwHiMD8YEUVKjlQ9r4ymasJxqBGP090Uv9K9AVBpJiCfECQ83bpaBzxU
L9DaHDqVBW29/U5WDH2uONx3ybE02HdQCAPB/v9pPuI+Mk+WNMotBh3LTaXN8cxSaPhRyuzajFgt
QBZnW6cdonD0UlpSP4SOeABv2ZNYscwF89CXx8ITrdpn0UI9Wbb17TFo0c7/QKIvXBTe5+QE1iE1
kJsjbQPicQC8fIniptBnPyYy8ALKLOfrGX69jaITLQBjTwb5j/+3YLJcJHBxpHz5eGgySdnEMr5w
590eJ7k/WKD27rgu2XaYY8a6FGqvY0p5QOElrbkVlVjJ7qrtzxaCoQHEpgJxqgwGWJJ8e9jKZ80c
qp1cYiK1PuDh4f1Z/uWwHuguxFQAdTZBbclQUSFlKorZAjGP1+89XRKM7p9juvLclz506OGvy6+x
BNsqiAvsfu1joQRXg7v2NmI3cG3SulAKqcsbIe9Kwvz/NPWyhsyOexUgBy0ZZOJa0scEhMOaM+yt
+6zV0Kyrp68HUomdscHxzjwYlDHcBf0XslFQIzYgB6/QgCRlKenvzLBZEv4pgKuo6bSIjdXIxW+f
XuT5BXsSuN++VY5ukpBBkattbQgDam7d+U4zWTIKZ14A9lb6NFb528eUQmwG5l6z1BAmcBCaLjEw
ABU0QaXmb3AypJ+4TTuZznzpRVcGJ9XJlRn6fq4kx6tV1XsAISHQe6gjHtOdSNcgA+vWcFLmFsWN
sq0yoLW/YxLYhk1fiZVSuCXpNVXKbRKpTqf7Vo0dpS+gtRPMdwJm5MG+gpk/7SFc5vb+vCBxu9iC
umElm3Wag/OQ21FA7BJu0t67haVomAAwd8R6uV3qjgLalLuMBl53u1x2XpTbp4Y0Sw6khbvAFGr6
0q7Y7++V0vVP9+g/Ql56NL6V9SvxYc4x6GXk+6gH2OgUFb+933yD4UJvppZBHi/Gkj615qy/csVH
eY/vQfPmL1c7oNYJeJw+EYNH6LNXb65jiP9DqJwSI6IO55Y0Acexxw69lvzHkzHWqjlEdRttJukA
+uviR6+kkupE/DWQL+V8jcZP5UMdJyhy3urycuPSqRaIc3R4KOUFHRQ7JvsKgda8CxEUucWDO1Lz
9QdmxZLIYaNUJIXn0tVOXBAInFTC3k2Lok3Mn/L+5jO0+DM3TzoaCUdqImiC8DW6keohmTI1ol1F
DOgmC7EgsA/fi9wlTTbHO1wFqlVTn9KYKyn2Zh8HBKK5EG5y/uOhNXcF/SMgZqs5/hS4TFk+bWeW
phxvZ/bDeeOoWd/LPxJEiA0WkvI7Pllv/UNU01r5kw+sUAJ6Xh/RVHCzn4SoplpeVqpfUjYtGsz/
BCsknZOMFB5P+2Ls4/85B7QIp3NNXQAO63VEQdTvaH0+8p2NKMRoKk7WMF9KSUMnVXuK8XoPNN7Z
apNVH9SinW9HQSKCsKNnRhNa6e+VVmWIQt1Qev96tmYqIcBt7c2LHxqAI+h6Jr6PO5N0LGcxrxPI
p1k1Sbuux+1XmRxl5mUnjhB9rjZzvX9W79/Z9jakk4+qfu7BY/OAZUllPRmjDq9z+gde4R8Dbsxa
S0cJU+ssM3qgZ+cVPVOYWadnxXyfsLFJWio7REx866cEc+MmNCZT0EWgW5EovjRzoSFz9DbQCNzF
o3lqWzoRS/Zl9mJa4cmMtaCWuTBXQgQGCrONvn89YTeFl4uc5GSrOyElQ6/c+KB0415f9qM7h6zC
OWueOl7zI1UezfZuKPzbzRoExAvhgyieFW0RclnePI2GKQp+4b+5VdRQDY8TQGAeOax71ndXOlRq
SlH+LKbb8iNpAaJq/WIjQf7xfjBo+uOE+kKDa3ozy8VdTjw7lQIoOBlE014J8tDSdwS+vkdtP23j
Pa3/ZHH1/XSUzho870C/PNvpy+1KLb/pEb+hGsBQsuvttFf15ya77578R46pbedLwKA6z3UezJCy
KH6tmQ+yEQaj+2jTQpEP4Md7Yf9ePk0BbwLU4O3eqXdxiRkVCABVOzDPSWBYZE6EfhGVO/qdpgqD
xsv2pl5fMJVsL+78jy4VFKSkrWUurcDJj8kGX1RF6P7LCWzb9SRPkD05l2rxEjkVDrMpASXocti8
QweTVmGAzngzMpnAfogOFY70wSCbnbV/GLqiqIELZSJqCE+cHdqbXCETdlWDbbe96JZ019W3DjV6
fdTwtdKWt083kwNdi3Z27o+1bk2ejCC+Q4E3PFKhwOf99YxnMtLcS+0BbpDmq48wv6WWUMXfyB11
lj4VdZykb/HkOR94yEQTtE/62bpaH/pcU1TU8KGlWU0bF1UrpAXqQAY3eHKuQLNrmBUSbMDois+K
MYy/y3hcbh+dpkFuk+o08gYoJmmE1dnM6nansGUhyNIipdMzC3uyAl5u9WVG7Zzp7rob++Gal55W
4a5kd0921YUDI6YYkHQIxVgT+8JNZMtiZfvzmxDJv7hHmF4SIJw6kfAXZPoaHAQdIt3mPTCF2sun
eSJOlYunjFKsq0hjhJUVgjpK1iFlmQQ+95kJ+GwPI/g2ZBeE6Id98SY3jSnAL2zvvV8AKqgAZj8/
KIEVr05MkfqblaJU4ZVDM6Ojy7Bt2uxTQhgc2/AH1kVlwmsGHA5L/iHwkfMexjwQ/rys94sNvRe1
qpO158/nHjvOrJfxfzQkQbdmGcb6oQWpUV/l+KGAEO+mmTbfWwVP1/obiwCnvMqf6ASda6lq2vgS
NdKufy6Wl5eVYcG+tByOVaxzOYEyRy3xLZ4tfmNc+51g2WxSdZV+60RRLfJY4Qx3mie/XrB46ACd
LXxZWXrg+8yyNq6V1jsC7KbUeRFZAjs4ZqqzD//jOM0/vOkjXpmwV7veFKiiERkJNgDf49uycyF/
mxksh6Uxbs/aJFqfEF2WMZBCNK3QCQJkTrgy1ik/7EvCEhXJB/2FKzcpyH214qkMZTHU3eeC6gru
js8BRioVn20qVBjgv1zKs+ZmCPmLtmJqPFBYChlUbkYYhF6wMkm7atS0y++GUKpzh2FIRH8HNq+d
9kFqDMDf+GPxWYVSqmqGZrc2ZGymz6hnRjIVO8qM4s4kt+3KQVJz9dYy/RzR4Ee1vWIOqOlxIZ9D
KGuX+QmAvdfXLoCCfuGLas4MSkY8v62LpcU5OxPeu+0zN4qI69DrwtScGo0XiVet4CLx0bbHwRNz
FecVzE822Beus8ZNnpISNS6WVHaAvjljvFmmPSEK5UbcndsGZIidHsM/ZZ1QZdkDniEVKnQIXUKJ
Ls9KUjl0rRk9QjySmtPOYDnpW02a1QcVt2YiA2AQ08epKNNxPUe+pPPSPS4EVQey0F3h/Lbxz/kI
hXU93/oQL3U0VgVZR9gs9ztp6wALy8gFqW7+gpXYorcmxp0OewzQzxg3fmESYrw5B1cXM1b8DINJ
iZSco0/cBU7rgfb8fL4JanbgAiabXn6DNfjLeS+D738kBBcAlBo24zYpgTFFB9Geo9yivz1dfJ1j
nJfRtKbZlO0AOuWnjcaeaDM3eI8UtXH/7YbyqEu5JujGUYWH/SNQOlmBZXRPoIslg/0lsrYBQ5Dr
tnYBXd2Loj3+LZ9aTYsXT5yyxxYYSJgqffIaQwzwD7kri6koUZ9leGoxOuA4or7/Yvxb8th/FNqH
B7bv8keSxIYko3sEbi48nm4l+5RIOznC6YfMMgw1twRB5l4RpfZ4HQzDWaSV4pIu3/iMnjKtBBXZ
6C7G68AEX91XyIshUhBxP3+Ch17j3hMVlvytem9+B9KmhZ0CGpUXc32TuygfGynGd6OU/cv2bzvU
PzYSkESzrlKLkfBQHXH9WiHmWbPxFeTRGj25mNV6kKlQsbs0fnjsgQ91WT5Ct1tC0zmmBRXz0PEa
g3bBPCGdBBhlPlVmwHgd5NJ3+V1ihe2zWbVQhol2ST0KyDxYgbvKeiv5Ck2nUYlc+MKAYWQzPdsR
gYbTkD5wgViO+jJ4SIFWwYQcWQu0YI6DaBaiQ84Ik4GCBbcLTY6ClhpguQ1Rzt5vbp93O0E2hhxJ
QUtRb2eUUim6E+vmxcEd0STPcz+n3vEjlQgbNvBjC1LGRnG+B8fv5oAN9tuWKg2L+sspandsREmO
674R7xbKJlX0aUzCMQTnqQZs9NHaaAfYeiEgPJc2toMOiJP1TseqvXnGm+8HaPrnxLquQxKXXsJX
CTd7UW7E46ILnUuhWndN1QB7k0GVWNwk4cZQMxia1cxUZ9DymQUa57CZir2cQ+CgB2xV2AtvU/hI
JVNTiw935CLOqp3OwdZxG32HKnQFKb7UBBMivDxa3Igfepl1ie2hPGvLJWIJD1h5fIDNQNdhfzM7
ZzGfG2x60dunLxSbXJt83kMAHjBWVc+oslS9/+MObXvcIqp94LKMwWRTNP7RIjAJLzQAytByQ4jp
dg+h0m6ABv7BemyRW4gyZf60BhgXGwFQ4makr75hHB5pzlM5hu4e/RAAf6aWVPg5Lz7USMoC966B
wxpq4RNiqEGHpXmdCpjPtchAmaD6HRDzO2Gxax6OwnAFXDCHyZhyRpQolYTTTyp5BcWnKOl8huhp
377gb4qtglv+JbOtrFBS8hY53uAm7/4Ejn9nSJi9HNYMVGjAPVsrCh6ckfMGKhj8YDj1xf+rGDJ0
VGJgMzRhcn7J1myb6dRmbEtJQBdaytx+J4LB2rxGTbX+wXI4V5mJOM/MhlQq+UOLYrr82jMz0T2D
n9j/MPN6ZsMyBL670LH1m+rnsSyvB8VZELYgD4mJFR2QzxY0nCm6t0kZHjHXPcALsJGqPvL1RKe8
GtcLzWUd4b8ROvSFc2FVQ2Q/u/uDiP2DTC+gScjc/Ocif7TqofKxNInUxoK+tdGSIEa+JRgY2Vpp
0d0YBdM2CzBAPVPcyU/0H4KacH9v4WE8G8/Xqt2tT0t3ZybBZxUVeWpJc+v2ew4kJ4nzC5RyT7Qc
KlhZXAjRgmiVwW5rPlfj3gpTZzPfmmmhlEdnhSgHv45OaM7gG/cHgw3V4hOh+CWfobTptsJySAfG
whkiZECbyeoMMQDXGBglgBJKY+tKcTaqLqL1JHDKOxpnsgLl+WESEud0jr322KLtcTjxWfTG/XUf
ziSO7x2U4Dt2qeuAimtlSK/Rt7wCv5Re6L8mbwtqqVI4KkSGiO8AyiW/PNGyJyeUsnZWieXbUlvk
LUyaj8bEjWC3rOVP9FZs9yKju123JOUD8au65KDy5NEnUaOcu9kByrZfFHXnON+bdAyJDtlgAbJY
dln91mPCPDHLl/9aqlwobc4LlDAClCMhrEG/Ex2z4LzPzg0h8HkyS7Fs8HPd0wdl7fGsw/9bX9E0
9cey+9ovj5F7fyrpMCWtWciXVSHHcqrelqALCd+VHTNqPr5InB9bMc2veKocTqOQZpYPH+XYrCQM
JYiFPdzV51+lo367/2T290xXR7a0Ii02+NP0f0gUlM9hZlCoPwkB5tlxS5PIfgFS0vKehMmx7AJt
nYs3Q67U9Xwrcd8gDSQYPZhIT1NezLC6hvfK33MoynwDopTdyRjQDim9x70yZvuogaVnWhFaxx1h
tQjRoponRyYE1oS8W9tM6Sr+wUJqHOazb44a0bSbP8zV5H27V3+J5Ezrw/662KpJe2MmHaz+daa4
MLz+LdU25gg92z6LM9XW9xDaNeEdtc1uQbuziWzeKyXuTGCXtJjUmGiFV3dhI8/JQP8Txtbivf1w
RmiisF2NNyJ8OAzoZp5XUOgl57ylOz0cfO5zS0VgK8DVOc31ymYzGl39ubEFJHOmpPkCGJMRA0hY
/3lhD+ManF2oJ6j+oTAptjql05PwlbOJ9Q9krRO4AAKDUlVGTwOIrdDs1zeM441RbtmlB4OqRAGs
0m/dg7h3juqsi1E36/Yq+86rkIyBty4AISCutlDh61eX3UrAx9iG8ILHH1/BsJsOQaxHZLjW75dB
MZhJQQScLRVyBCjEcmxaaD1n1V9PHTr2elqjwfbDyPhviCbpYzIn+N87ZAUvkOV5ubO5AL9P63DT
BwNMazHv8VTPTI8q8vbnvsDVviiuO7rZ1eTDhFDLUfTKxRBJkxytZ4pb/dl8xvep+qdt9qRyR9OH
ZOszEoOYaUJVkX0AO91pjgpM/yG7bNj4AK36fwdW1GTeVEDm7BgrKt7iFmiuVa+OiN1/ZEEJtTbp
ktTPdDxdb7rClSB7RsjPo9Jf+q9PyDLGe3pf3VF3ESwEtWMMwdnveWK1Kub4qt2PoPSP980GGbzZ
eqFCB7YCG0NUcVBkZE3fUx83Y8zvcj3g7z36LGlJv7ZH9gDfKzfywIQ/JwS5/HVrgQfpiJ8nu5EM
d+QfoEiu2Zdq7CyqxOCneSHwlDxGE/Ts2wrYR9aGhwhF9pWcd8iCzieTNzhnE1JxY5AYzRU1/BkL
zATaHq19gsUa23b3knKhAOYHweD/TXQ3ICybU/WsUtB2GOxb0Y6LcxjjIcUFTf/JSZ5NZZwKbg4t
DRlrS2OKojm7TeciCWazOSFVgusfRQyuSvoXIzMt6I0ibqBe+oq5IKPmL0hgYCJcz1YYXYy1GdMP
qpS0P4ubsiHnJMy0o9g1sROWfaOW5covjgF9O92yLBVjTuTRIQL4P5ttifmlycvBvQuTi5+a4U+d
ksn5hYUGGMmYLKj0cZdjGQhVVvbafRRl0+VdC1WTYvDuceEXoobb7UPpodpPokPhXbc9kmPR4cqE
qIFmFEU4Xb2p7++Lbtyc7qZew0JX2EpL5Poi1TiZG7zakPYkZ011DC0r2rIbchrwTl3bvqJauT/K
cLo3aPVxoR8CMrew8azJ3UWKTZjcxMd5QNCIKYFeyMbagQQrN67G7yAiOOKW62anTSvNJB4SYuYo
r4mFi56ITkp82JBKs1/DdupjllpvEvmlfYcIYBaeANXOPw9xl9L7RJJqTawFqGfHH5/galzMl5H7
vSY0+jsDHwoeeHNTNLiXhLfjQA7d7dcvAQo3shO7HT+Zr95yLJ1huEoN78Y/frbE+UzJrdPWGSBl
TeFMt0fGbzKPGbNKSXktZ2VsUwt07mqKvoj1FJVjv9TFMyEDR9K29qQdpE6nPKWo3a8d+oVbLCmp
N6SXM0MKu5R3wcqgtyB+VlPGZBgYUvXJOY2rdxqPHxCI8Oeq8xb6hXHdv2OBsBQrYUsEhTLQ7M9W
1LnCD09vdb1tYL8VFybxKZwaDFMc8hHrytmujWa64saFfkvWoZUCRffl8fRJRl0sHxqFDuzWun0e
5SjT4KDGT+pEHpbZsGsheSTrfvCu5gQ1UjW49GR/9uR3Ud3ioBffeHtZgPCE+iyC4ox7FTx77rbP
FF6B0fm5SbkC6aVQ+7OgDW5k7b7GAOoYAY42rnENgrfK6oktdlPJL78geL553mqVQav3e3kwYc/s
nanz6w8ZcUNKWS3rkb9ydLsbNi6c1iJQ+zfIRsUDrpgWmHxAr8eqv6CoDDz5Czcd4RIgMQDD7yyt
9CTdZXPpmU3iYDbjeH+tlPV2kkP1VSpJzgDhmPbCBgqFmhEpXeDTH1xsm1hNDp0yC4ax0FvqF1NF
AdZoy+N0beka3IC9GSP1mWcOiOBm7EJpI27+ssjq1/Ba5iBqLX7Sg2woN8tNQYW/iYe+U6epLjjm
q9dDGAQErwkr23KxcPAr9wiIQgYO910vWieJelM5GL5Lnnzl6Zhf8Zd26CyxZd6XUuW6AmTzFD8y
xF89N11fqimCqZYOSv87nn7aV7YnSWnVxquRGsc3JsMj0JJ46s6tgNp85g3AZ6TL3PZdYnbNlp2V
+whUTrMGp+8dmK9QFvh0dMyxigAEt8Wc/ScHjVfvlWevBKs+9cS4ohSnvMxoULRk85M21PPAdhYJ
aCimpsjiwMHEWoVZtC3II1NvAJbsAdq3e1/Xxg/NIU9JHN03uHglOex1MR1FWjLpoEA4LtDQ9GJM
vGDf0QbGqXK07CsG1r6aoe4w0urWjUokdlIQMEf9zKwWzUf4H1+HEoqtwxcalU0q561HrYo9MTPU
I9EE6mf7rGxtUPQZMOwE0yHCzJSBUFgMexJWbRvzfx5Fp1vVyKP8/2YltG0dBdAemkB4KydqITgl
spjNpwQwi9oiVB7EmBviFAE5x9tfkOss9t81QL6JAniu9xGnedmEzK4VpXbQts0hERFzI+5Yt5nk
jLY987zM6aptB1783QMWasikuebDc5pUfvIxB3X+TO9HLqPzIAObwX0lEl07Dx7XE/HGTmNFBc5a
vsGrAw4WSDdePEiEYuW2sYccsbN+MHruFBD54hV+Xd+jow84p8a6NpxyE/sHVHmonI3A883w7FJ2
7xV4zDSp66OkG1S0OrUuq2zZSIXneP/4aDCfFVWpbwKKrpUkojJjxLEOd9S1AjQMb6cAKvgMm/hr
deFoYxow0k87rhCxNw3aI9cQc13i8n8oCvtdLfvhoB//XOGr5tVeEml6X3S9kUL/jO2lZBR5qNbT
ZXb/YKrWMP9kJLTa6R0TnBBfwj7zBnyEX4FwzeUBuJ6l2Uq5h3Py0WbuGw4YtwOEmIxU1zdZD5Dk
LaymPqC12qJ67XTy8GaQxuqg2syMupneqLm3LEWjIqS3cA6RUlKj+Nj88OLffMCorW1OLDuQnVFi
Oo/0n/CzwCAXQBZkO6Q97u6uVQAWRsqzaioa0EusfxYnuVcc7Mi6ZleIKw7z5hBucB8dg4fyw8Tz
SngiTmC/h93L7l+om3JYUVgzKPaVR0xuZKJsF6FToed8M4nr0HqVZ2zfG26OlyYdb7BZfoW2zS0C
jFNt2GBwLDgUtxhV1RzsFT1dt4cyFf9RATDDD47yW1LH4S4+HRm7m+CwPI1dq6Vel6NQhbGISSsO
IzGMxPL38XddRPRHhSNBHCKsDYR6zOFdQmOLXXKkesNh/O+Ht5xqHl1PM2727VbUXgns2Ki2od4c
/pNc7qAPhFxYWchl+otzou2ZzC1jZZL0CVMfGX4uDOcV0IdlMoQOsm2hyJWtj/AZmXI53A5v54z7
fpZZdpCmmXvb0K77CSBBqbujcy5J1hnwWfz4bIljqsX1cG8fTcdGSlDMBDc1a7ntOKXoEtv4rFNs
T8rYMjrmgbji8lw/m6tSZMfLXl1TdmX9yn6Ht6QeakZi6RGUHdrXWZbSAG6TvCbvLSzx1aK1OUsY
Er12+AC2WkAqyxXYuPI42xdbOQdnmroLLP8ZyvcqtAo+WZLOsFq+Iah28zHBkmnOdPy8wBaPZVEB
+sIpXyZuZe2mI4/GxUQqJa/2hxp1USfjJvxlC158sCe/itMPxHna2kqN/WFbQ39XdkfmnLIUL2AR
bceFpL+j0OFskj0RVpN9iofZyZ6uVrtlciQOo0ZJ0HBrtfkSsJ0d0tsK53mLFPO6D57YvDQhO15R
g9Cf1gyaSUEzm6JAEcIzf/8oFzKP92U4DQCMgx43CuMQWUBchxyIWkv6/2JGLs75ZqaKUwThaG2t
uY1z0ua2hilQt0Po8VerNwnvdh0yTxcjgsh3eHooV0kfByMtK92uww2km5SkYmvOmUXEe65zLFam
igpnKl+eTd0zBk1QL42qSKHNMZeYuoqF7bvj8xwno+q+l8YttmPHKkfxHteR7liKvor9Tsz3EnzH
jfACMYemaGDV9/j4dd3orEpybR/ECYXHvXLlt8sTa3Pq3Lloo726aAO++GPFFQvE0OPuQ8T5dtts
ksq1NP6c9tCSIfBCkItYmV+jnXwHIy+YIrhCSpSdUReZeQqa+uCD08K4wx/SRJtpzNmvKGqSG3+7
a7c3m0HDkpCobAremDw3+Ul+MCJd9uEhWPgZjh2yDtnirqoFxY9ovvycck5hKyT6f0Av+5VhYy8s
3VASjbMd/u6agW6/fp5HtFLokbcdoBCCgNRft0KIwvBHSb4rJTgbt4hvEHDL46l6mb9i1CuHDztK
F40DxdlINd/uA4XJgIbBQHmkp8JOluqHGVbzi9zt40ojAS3D41p2Hq12DXkJKm4wxMmAmdxTy9FN
PpWtLl58GipJl2k2edOX3cfXztO9YUIi98TUTDrEcsAC4VTvlEQa66AC8xt5vYR4vYp/Sogh1W2k
6hPL9YihU44QaWbs2sgksk4v0HkxkcIQJYRjFjedHoMUJibjG4e+abrwDlclJlGw8ho5ESx0yXk0
39dfn9IgvZn0RyvIqEMEYYwthWmhefv0f7gsoLImfqRJy44NqjBNjeAVmRJX9g6YknhZ4NzgJ2xY
/6X91R5Cl7kxZ4UuMsS+rRBnNusuBw5uLlLLhPwGMfTkI76mxiyqALAz4oyYHHRx0tBz8b5FvNq4
+S4Hw/qk5i/I/jkXswytztIa2AIf7/oBpMJN7CIIpOZnzVtgnYA033ytvNy9CcblIxYKs0gCpuIW
VPHk9Ya1bzqczQbkgVA4w/I2pB4cejdnSE00/vwPHLawAbnWBtAfKsDqPAky3KOfPOThRrqLKbv0
vwfDbVeiLIXG5U6+HU+YYj7tMyCz8oBwFjhoXt8efCiLvg61q+lxI4QWwuquKqUDO5xANwRw14f1
cvKmMY/8CuvPiNtZuURQYZMUc9Vxhp0XfDLwMGZHcj5TY2hzgWHoDFQ+pImWxFbH9vVZxcj1BRTr
V3+jdChZSDoqaDkoTZrRUxoBkUPSPTPspmKVP6BcFaGgAa5Wk2BsVj92UauZjthcSLrEU6/pNnAN
S9od/7CGx/11suLuz3uNYmiV1IwEdT++rEzv7Lc1lKXxwQ/U4I+THFbCU1oNaagIKtsWdBSmUm7t
7DKRf8SgtVS1Tqa+DuR3nmN3nIVnDl/XGbgaxCO0yPvddKrsVWEqzwn1u8343VD6Hv/B/Bp5bWbF
m5NH6U+EjotkWVDiCyWzs/6YepYdwY5Ccr2mX2wHq4h/RhzSOGmQ7WFg76Vk2+zB/nFXbXkwYSxR
aEKtVdfcQDRNHD7uROvDQ7k5chFFXP8Zn3Vfe0uk/mrvgjb5opUwae0q2U133j0KPXmtDcIwYUad
EW/fTJm3HKUJCtegy9CLRHuD2mosMsUhz+iB9sKN5JgAH32+QbqKh7VdtwXPB5DRO5CeNXEpu3So
6shjeksAX4Wo7qIk0WVgHvvp+GpWh3YZBRobP3MVN8J7FlbkbDJaGPJemxQENTTYbx/x54f6ywuQ
UckGnxB9wqEwPEaQ9W5DhvBpIUfOH0qDPkkPviDpyyKtVLpWuwFqYfNoa1XXyE0erkNURwHr89KU
Ufp+xNEYS9p04y+uKGeSPhYbHodjOxP6k0jAU9mhEnG0KESik3cvCbpW0yUlE3FiEEGZcsHybqD5
QlujeO0ig4zYa4XLg+OiDCs/6osV/my0Cwosefw4KRKHXDL1BMQysd9k61JAmk6mqBe1wjEHaLX1
3I7M9MWZEScaDCBtxWs+sGIeEeRQSfNAKxZL0NPrwarMGa0jsleMAaWAkSAk8xVlXsOH4+WvSGdO
Ua083vO1owTchzEp6AMQ47elOQgnF5/SyHveHDaxxyQjN4l1Z5tZQ7OjKFheZdXTHW8bkPBQ/yWx
neKnjJ1ISXLnXUFWGeDFWomUM2/RL9lD7t+7pvmiZi/y10YQ58/ndAPBpq4Uu1xur5ExjD6NeTkW
GkNLSv2MjPKDfYwT8HRuUoNqOFh775IjI+3rfQi+gLp49DjQ4GzXiAodliZPm8USS4F2z1s/cpCy
mePvsM0wwRdXKYZ+7PSuX0YmylmF0j906BIlVGomh7ct6xuTezsTX/MGcHOyanJgAHveLcfzsJJb
4w3b4r/1BwUMjDbNNPecEUzz91BO/GP4B2jXovU/7KP7SUmeHUF0snrfaPPq4rxjmpiXskqmJCw8
bQ/SVd2zn4EFFGpZlSEllPlQo3oTLCXYdimsQ6QM/jn6nrCOgKu8TWV7rSzn4rwIYKEicBw1l425
kBY/W/NTrq/XYIiB7+GYx3OzvaM+Lwr8a3KeQ2B+BXF6fae/KNRMw0Fo2uqTmndK/PyNWf+uwy/r
iLl6A25oyr1Lc4+xmEY6lcdrMj5Fz6j7Mo9ChPYeiN6We5eKKcoW3y4P9oPTGrapnOWDSSQGFJU6
GtjYQFbmWuRtKoojC+K/3dMeWFGBKPM7rcwxbQS3Ibwb+XiJ8R1MD0U7oa3BpKun/dZ9tT0sNtjP
hQaHkCG3Snjx5q/GXFJbfhOmGwDSE+YDiAq1oZ1m+o6VC2IZpb0McucexSpoKppgM2sYBYkCYEk1
+83f3kc9JIwMgc+pdYQLOX/hxX8JYqKjum96zPUa32wNVWEBIBe5cbHuYcq+KMinsCJ70h6GmeGd
3QihbFuuP04J1KehsWQgKgOCPgx+sclgD6YeohdJhmzfnSJK1LnnYkoYW0BMm0+GZ3fhmN+l+7FN
1BBF3WjbFs19U7B8STpTfLAM775c/bbfJIQu3ybiF4fe3uMZ7Ys4KGECNqZnMl2UVT2TRxKkEnVo
1SsW4oyws5eI/rL9Dm1CSCQffrNnid/OieG70MHwS1GHJG+yfhTfP0ev4T2JsvYYw0MZBWDpCJDA
MrihtZilNuIpL6VzQaGysah0b/HB7joRfGWF0T6H1z9KmRPnWTKYD4gwf6017S6+PWG1u0LlFDA5
okbkUntGHDxQd1ZHrccbldHMLnn2UrN0NW9PO0CiD0har78hne3LTgnG0nHK8K7IPbXlUP7gcmkc
NryeX4UHoMoU/QO0Gjv4ksddE4xXuPqqk/WvBafb+ZR6pctMycMALcUzJubXcPfPK7N0eH1Ch2PZ
7tCbcnBuShJ22t0PhRGRHsMLfMemMVEfPZJW8epnZMztY+xqhcMXNSiwES8nu/75w+U3Xhyff2kw
HzFsT4IJCQ2YSXS1L9HKJhPPA4lYmaVJiyar3IlIwnJtjRTr7zARRS5Qn0qX3LAJwVV7og5OIUDn
Zay9wNym+h9JnR7BcK6eARCTo65/kLlz4TqRgAMngOnRg6K1CsS5PCTsXJvU0hwMeX3lD8w5jH+Z
7y4o8dgHcYM0bzReAWfhjv2U55oEqsZPWluwnTAKEqQn8TdJgRtXJAG2va9iWmB66lyIkv+65NJ1
MluqDUJEfCYe0j0/Q1M4c7AhbvXjpQxzIKEXoneOw3rNsWf8x+QUZK6Xh1a+0/rRf96+JzhWykE0
hPkFRjZFgK29CKWckdOC7o89VaCErxea+q2ONZokLtieajYKw8BocpCUziJqGiMUi7Y859d2lrQ/
mUEUI6NTv/K2XMeHcJD5NfYUXhbCkNM3PL++LBQm1GxTvAjLdP+B92EXZDnDMSidThwuPqKd+h7q
m1Kjcxo8TzUJ4oSkl5kRLzFRWWV+s/mqO8U8yea3Rp1tNH13hFpSsxB7zT3xyWyLLhn73b7+pzBV
W6Qm3g1upHrmNZ3aSjlzWaC2t5X+LxquGxYka3KInESb71BW9kKdVQ2b4LxpVqZWmIdtQwq771IL
bdhVsFpBrgjHSzYvPsHBpZOQWDEi0XuWYAwLeu2XL7tDLAcb1jdKQuJtSFidVSQX4vH+ix5NpgPH
L2QlwoboBBpoRtJltr99k3DepBS/d9SfvhGXjPICVWCUtLhELrDZUR5/aHCcl8KlrNYpwFwQzFCX
0m6mKhrhggTNQXMZ0egJOZrzNafr2wlJT4cO5itjXGaJGjEpbbePcK6Hrm3NEhOXLTToZbWXqD3P
xo1tsnPtqewY6KbKmJzkEuMOyAntJ5NhvpE1BgjMQFgmd7lCjrl0T5BA/y57noD5TODI+t7atMoh
FCn06S8FMz6vCd/t8HmIcD/SQbvyH7RJ15AMJaGri0s8JWu7OMOHkVykeOlAenAR++eNrcE7QFaI
yHv7lRTlR4RasSMgUHogjquCyCSM9n9FluQX9FTw2WZhsBQsIq23XNWg3HmMTN2QK3Ch10IznTXW
wVK08tg/aGYS2MzFcyW9BsHx1Gcm5jnoovIp5R8Y6uMfkc68YH3YGvVunKwl93GczLkPiHQwJ2Oo
xclvM/WTBcjmyub+g1Xsn93hlp6AucnyshPZxj4YSAyCq5svMzPWSVc5hrNwtwklu23C4evkGE4B
6iTlQWiqA4gHGSevsGdBp7XaFjE4U9qda/cAnUHADIQKT8e/PRlR6JMjdKkyzFlTdCTqHHiO/JiP
wLzFobhAMuQAt/sJieibTEnk04jkxOlm+bvYFbTxDX2VHEGaijv+b5vtL/i5mnmcH0BAfgFwWZY2
6jCoBQYOR7MhURxwrOIuErhU1LNboLqHFWWWl/198kkTrOpUWMmvITe6B1A5mBEpylOiDz7o0pad
i28yUjOvHT7PzNplmVfUwDhJdefsI4zuUacRZB4EhGXU9/6R3UeAG81bE65U91/dZbQorOgFzTF7
kfMJe1J8TvWh2udROIRvn806iEC/LXEkN10kST0W3wMzHeTeHH/9KmKPv5hZJjZJNBOseRnfEXwc
gAfJ7OXlrAiXrT8R8g00zDodsUel4GcwWs+RAFlIyuYrVu6eo1fUyFcW1IAVds+TPQzhy9QAAHlK
6WrsrmUurrOhNAGDLV8sueA3eSckrc5cBpYMm6jkU0aCxPTFwQHavkyAtVreDQqb06WOKi3hztCw
Yric0lL6zcgkzJGkKdCLhU6yPx5DYmHT5Ds4l84yBTVcQT6X9UpXWwFmnkUm8RGOWHZNA/5flAo1
6L9iBTOWHUgVwQqbZiGk9lsVNi5lca6tjNgOiyY+9A+LECaYdS764kcB9OjU6bhvghrkCCSeqV7z
O2KoN7W8z59geflQhKfzzscVz2m1gAsZ9L3ppH/Eyyy8WxVLHc3YXLQQLkIIbf2Ne5EveiaERHJb
UwcvvczY6keR4bGIBFxgk5IDwxSvNw2SSSYsYUOl81fZa09CvpLqTf6Iu7lB9uTeJUOgz9Dae5Nh
V/a+BObSX4GtxUtNRqfEXpn2T634N5yaIW8IjCUCuzI3knP0L0WMQ+RpF3QGT+rX3sDAzEFAfKHx
jCcpaD+5dsdgOfgQ2ECsRQauIhxQy/SZBv367/1TcelcWVYh5pGvF1WVjDMUwfQ/CVuwT8NWAUze
/QJ8g9ptXOj+ewhKf46YPAUZQqLpBYhRhWzyHHEZNwDISY66/WLCQMlk58+9l9ffnwGGgWWCb/bP
wfPHBya9U/V+Fl5JB0FQYK+oLBRWXxxSyNQCak/Bb0P7A4VGsDL50+PDzHW+E0dMoPXd2ykqxU6i
Qvm7KmI/UUG/PMi5sdrchxXO80SXvOmJW4V5uBQVZ+3SU0Vop8EKbA0I78TKt8/UK1rFtqTKCn30
idul9DSvJZK8WiCsY1kDA2290UZoNIzrBppU19SJx8u3uAgix5M7ToDYSLR5gF6+cvCjchpWI+g5
30uIMZmSoF0alfaob88nAVh8bygT6Nkqzwzom+VhF78J2gZeQY+quRkDeQkGMrZ1gWgaJFZRmmMr
zPF8wLOtImXNiqFhoWvFiPltXlWDx1pjOvAbDZXfGHhal8C5UB590gDJzqIz2D9LCYOKJmS+76ic
84BmRb4p82oAvbHXssVUgT+SP/OC/xdOp1oPZglLp3rB6jqWZt6vLQae5Y6gpK3UrZGyXSKiv2xh
tkIwdc3lgBDnl2oPvtOiqyJdEEqP9AwiU8ImCiTsFmfDhVe7HjPSuLKLr3D6dAoYVDfNoCRGq8lk
OIIDUVEQHzuxMhsLaG3yMPMKMSaXoHHcV4/lQqwsiH4R28c7PRK4E1eMHDVgcEBdvAz0BxlWgDVb
74ix/5p1tUmVGgeu5loLyTCzQsOcDoAZHcuY2G9VGs+8oOzpABZURvQqlLPGfUmOPotmeKisBoGo
JmfvczkoARm4snKzvyjcr5G5UosHaFURbvJOdBQWFLlogEjWfEmtzityRr2mgiZlT7kZI4ziwvol
wIakAFyljXFMH/axdQu0NjwWRk59o9yHQHYiFoTlRm4diOcVLF9ssh7rrvdrMoDSvVyrZkqyA1Gg
URyPMz1bTe4ixgbpLA3AiN/zTl+9ZYTb7c4fXbU3FF5BtjLVmwCXo2pxFnY7OPlgtSJfJMHPzcyN
nQMRln//3oOXjokRuST5+d5PRzb5L3p6JpXkfIl06jw/U/kPAqvkP0RqjxHniFTYaLUKGQqdT8Sc
tV/3oTBeHDdfV+K0n4yIj5voJC8Opkweioo/dv+oOUy41B9CejUOrYt1N7I65X9IK/MiDhXXcHBV
mEblTEUSWI2WgyokemdvnbZYChDK8UcCtuiUZPdT/P1Vx2s+MzM5TFGxl+U2IdhnmEZtUTfk6Ku8
BtX6KzST0i3T46Gr3UuSLlv5RNGo7RqZ4QyAq99Avrcm9b5f9E58Hy5zf8R9QJFfHoNdsUX/m4r/
EuRW7HEzTi1XPieeMWUQpXsra05TRQSqZKZbHG+TLkRo8qgrXWAnyihAUOPqbNAcmI3l9ZMDmT+q
bwztB2YduCTW/b/ecDEJblzgXZM+QQGPxgOoGucS7pYVE1XcqFvrTyDYl756Fr8OxtPxd4zKrhGc
38ZM2v3uq/pjF9hDE2yitMZCA9bilXV7o8vRwUS0Kh11m7mElOPTqhAph7APBvt0QOSImvF0VF0J
WKbp2Qdk5B1gqB8jfzrxxMorAoO8dBIegTNYqLEUsRDYBV+h14QakyxgbY1nN/gNPQvioKzyQt/q
hxq9i9ulhcZDBAMAFMMeluyxm9Zv5YK9xRlFVNDEXuSKsuncubUSw2IwnUUvWXh2v6q6u5R6Uh9E
EBr7NBGy0I97RYoAD8aHVIRWT9l8I8YRcIUxgnfsva5rm47bhozXbgElaFFIepDlLwUz4UVlqX0p
/QeUdeFyJHsmYNv+V3YHegFfv+ahU7fglBBqudcy/IinT6p48eumkty6HFOZOLF+Hdt3+THDFAdt
ohYXipHbJqizXg+KA6XJAmnB2DjGJrNFwqi2V2jEWSLk7skDUovqxNo3tya+09+MkypHN70rwySi
J9tBL5Vs8NmRgHxOaq4w3c3SA6X4AFddE+1T18UNAVvwqs6USPYzyZjgFUc0LV3WH6y5kqZWUjWe
+P7R15HFDSjucvjIONgHY3Gd/TP/YHeXdOUGHXzFeIIWiGfpgg23D5lA0/cL1viYPon1+9i6SwQN
Pnc1rPHCVeFfIy7kujQqT6TBlu6MsPdwX2qVLooy1pCorSBP1/XsLSaHfJUzKAt7Vn1snb56lgDX
irfjLGtO5zoNb6+zVZ7v8VVVH9H/nbnFoyIyx7Diy2WMsU89bkx0Kr1hPQbRC/eWfnJ9+u1o0Juy
9HO4bApWwhCU53T6c5mWwZqRCh/kRZtB77ErHKAWKRltLlY7n8aNJgFAbS8S0NwGW2uFapGNTysR
nFcAQ4akxCOCA6kf24q1xQzzGYKDT7N0AxEAAkzMCgddOpK28I3+yr/+mP6ilxzPv4mGUOEEl+wr
mNQ1tuQMBz1xy3i7U17TS2UWS5AUWctUw5Da04RYvJZMdLocrlIzfT3K1XtQvK2IZoBL4KCIKEwI
auM/q3DrDFEADTljHfeTNqo3IzRCIGG1WEO6c6bdP5aOalBItguBGwy2r87lve3Aw7pRnf8GQefz
ONgNJnMz7OL7+KwH7Hf9v1IUpFJ35VsyNHcrzBVlt39rz/0602KCgkltTWfp6bcDeII0T3+/Q0cj
qSfTUgd1qzGa5Gy6xckZogT1r92Epy0AYE7/qAt6ElItDRRrtL+eV6p68PZhSjrOFd5fQKOQzGaI
8DONH391K8/R2kd1YE7pqaVD1JHcfre9XZ6cdql5tzFe8cKJwtfQ3/olefOGnr27g4BEP3RfDVoc
TS3kr3RAEtbcpvIjppdjrOHNwB9DjVZALjSXkZvANTBFVzAmnw63mh234tfU80ez4lUODmIh6rE+
Hhl7GG5jR5PCse+R7xJz6er9zxya8iXcAbJjL0yADnMs5W5oBjRUYIIv4EhCn53rMs+OkkgO7NKL
46kDuWDX6ZKcOv6mKHMNAOgy/TA0lbOWx0v0K5FdNix7e+RJ/iA564BpixKpo6reKwTcKxp4mREk
e4e1E/54OZv74y0XIYtfR+Q3Bx9+yt11DSW3w83gGNA86+bap7uvVo69MxueYEzKZbVHIEw+8Ubn
vQFKZk4ULtzPCovKSeRj00rSCQddl2kVzbnhRuVuuhZOKKPGv23ieWPQFsWyXU1aDHuHB5rc4+l7
XdI+DbxcfVTnQSQ0sZ4c/oD1DX/7SCTpIfqJwN+qz03kFz65g5Ga4yCYFBt8lMz4qAo+Uzgf/nrY
OdaXcTrOG/gXdXPbPUZjSUKaw2J6NbIsdh2iM0OS6BPcmueZK46HBKhlG6ks+XcKvDTlu+ututAW
STeBo1h6g3/cb+5RLgSmIatLN6krodkdFlOng+Prbk/BLPiV0NPzF77N9GYwiIYe6Sjwq1bXKb5P
rTTuiJpEjyJuHBsRBxmijU80j3JSXOAQFUVaTaKJA6+abCZ1DcdInrBAr3jTmLiYjWbBuIey6Q5w
jGPavs098GBRXxZM0THhNL5MvBtwd8bUC5ZRjAL0yIAkDjCGffmCTVTJMws72/3PVG7+GwZgwaDw
dQsHUJteflMR5RZ+DNqEii5hrNeIjFkChdHGRS73FRDinyKsi/ZlGS7IW8J0I5PQVJeBPZpAOlFk
dMLtmbp7M2JekdQ8Ww8sBWxIcFgPDa6rzRExb5EwN7P+CWXqTa98xpW4DtBJFPU7vs9ZI0JjvbL6
p+pBPmgGyXrAwCJyk9ttG6had3OdGBwKUW80+HlXXqW5tJxzCATJK3BihcAkGgVMkOx6Opn4JrZb
MlqXpQmBzsw9V4KSq3rP7Y+PCoyJ38us2LvYKLhoxcAko/t+jhBR+tamPBa1dpKPwZ09N1rdzeEK
4uMmxGVTtvqec4AFMetvSSQ5DYwv9TiziNMcKN8+JcV5iYMNDRPLXttveNx9Rz+71m+OMkgvsbPN
5VuEJ3ZUzd2B+N6fQbV47qqcNhRQp03WZzBWQTVqp4mG59HNz3Ep5iae1D8yWmI8PjNkPrPgiqQR
5HsNv7f0hBG6zgHua5XpXMGUVE3a801+7spI/5z8sfIQ0Z7dizX3wG8kIivh6THmVkqUA5ZFc9ni
NTkTpnZC5C/jnDcA1U8Td7gNdhVo/cl4YpKMn6HmX5T6r4KhO+iHCBCQF96435atV8OczRTiwMXc
qJ60QxgW7WQcBv8p96gKeEZ6e7EvYjFf/BcVzNPXqKInTN1sH6jLOjMBMLUqLBKahM+I3MQlifJ8
34CA+esIsas/5R6yEpu99PuigME7A/2MaUfj6mzQ+fVLbWqt+oVkFHOJEVn3bilVV4K4KMVGUjKg
mDFBTQFZqCnDceugGQQdFBMUr7NlpdyCeqiAaloqy78vuyf5CNMois59OtMlvN8ftCev7p6Q7nps
rWGihCtxoHgl56e+7pfUOoTqNXqvPRQ8IPhs2E35y7HnKjRTQ6TkNmJBgbHRQ/h31KiJDDqcSetR
s+FvM28R0gpAz5gc105OJ2nCZehjMDXRtNxTwHVp3TeOxph684lZT7L0ZU8+qylNDl7RhQkHHu+B
lPTzMO9e1XsQJIMA/FYAhyHOdKhkKogRnxSK9+wU/i64DEwVY1NWoV77H+G8PxbIPpxqYPCZTD5X
81QYs/czG3liXsppw1AmYvnCNfCJ3+WUQ2ZUGirj2JnnnFfQKCSWuUH3nc58kEs9hdn7Xbl1chAL
40yGFlr1M+zM7PHmYQ5tST7/zQG46dxVaNmOWXzQiIIK9+BjV+qbVEE56XIrE/2YfFQHs5I3+umo
Qs03i/3XyTK1HjjZXE7nIRPxgy4S2gMKeWjk/MoP+rur0ujEciwMNeT/m/+XLMAfbteQeCj3eojj
VL/vK+1chI3CzDP0Q8f6QvrQH3mF3//bBdvOF7eCBxBC0wNzlpib6jOewHmhgTGW/wPVI7hZO5bH
Q9rX7Y0l1kBnlIjXQFulKjceJGxWf//jeqNyo+lTuCTPzln9cSfGmTBLfOeDTDcFGD60y/7qg4vP
paNOC/T/7k21kXqU7glqwwPCDwJqnq3RGOkB9ANFWkdcRnE4LDmeWU0f/Ep6HuzMTOG5i2j72KP0
MdZVN5Mu4lftoULZWdUP5maT7rgkfK6jhm98UJgpgkudz2dn109QHV2rCeYtWr/LNJTV4Frrs+Nk
nSeAxOfhm7UP2SahUWcvvaWTWg73+hyGkIHwev2O6L5zP5m2+fyrXbq3XIoFOPqWSzxqQP0QAO1M
PCy6jjAjuElZxk/zEQme9+kdlM9fas0uwoW/nk2jR4A27aHZNJnUv/zKjAli7ZhDCyFAiPqsoPvM
LflUDNcrIsb7iX1H3C6JFVI/fCUkbVrU0djW+DZ3QNvILztWHTaRQ3OwX+rM75zzQx8GLeMMjOOy
QG0D2TDnEXeblvmQE5jFKuPlt/aUYapCaxwzuzpQrLukrffyZhBeMQKLZoYE3HqBJWaaqzdSC/QE
XIowGLyQcOgEyNImUEaQFdFcNRzLBwCLX41dUuH2CarQyrliYRMwLm5crMHJvWOvQ1wdstM2C5BI
hqmZ0X9Gfa/sZNF1VzsgVFAWBCd+SQl6OSn4UX81S/zvVLvqDG/B5dlUSEWWLWkte/n18V8u0u4S
OZDfrgczR8MWt3PZ4r18N7OCFUmeb/VqczLShRe66hmSXpHLvX1IdckosoX0rn6DKsfxwrzCbieG
NgCjkAF3E9pUIahXScCceaHErYIVBGIXGzUhciIgDoGpQ/6CqQqm1G+VNpSSs/nlxv9kiaWFlUa/
YH5dzMJliNniHEAi4G5a8EOum1XSxpDEHwZf9BwRuhPk3K/zUkoK6VU0o06eBEVkUKQN/aV1TMTV
SZZVfYCdnsm4OzLjwlD0AN/ub8shLgVk6ALe591yjQ/KmW/DD2+tmjIdMcit09Fzd0KlHgCxzhOH
wtsdOAOZ/SUS0EIdlTvZQq9S0WRJLrb348/PLw8D0KlFnArBgSValrQWUPZz5/l4h13LH00BT6E1
GWqevyrGkh4UKoF8Jed76arx7jcaL3Gc/7C2GpMd/naGQ1mqvm+WyDVc/BwBuvSwP/EeEVSr9yVF
F/Hc3L0Ogf7w+lrHJ4SJL+0om1P7wFogBVv50KXS315rPeh48o3p0+9RnXYX4qVPUDVRHG9bdpSu
4slfXNxRhsur2wxZUM53nLA9i8aGXAoS5IyWC9t/rVcdGNlTm3rF/XzQ5bTW4qez+ZnULTO0GwA9
s6TVCY4dRIheRC2yoBeIhQuikuY+TQJGi9XICRcK0rzQWGLil2HBdNBDGWArqP9xCApOhHziN/ud
ElbgsPC5bXGt4LAAJN5dN9G16zXtS4um109rFdgGOuQnXlcthHWZWLoFBND5R5Xd3eiWaB4N2yB6
aOrP6gywwJCEAmJN9s8hHKbBcOC7hV96moR/jTg7C8CNKgtYOBGCNeVuQ0GCQMM3n86lMWFlrECI
4Ni3CF9FONU4pNABaVkmndeoD6L+N1cIa6TQWwiTHHve8lJnhlNL4/n7cuRvmI607eQ46T9E/P9J
abtjdQxJ23nwfbFsnf0bpc8ThoENNOiAKUcPClQSjD3+/qjCPxMPuUrPUWrJOhhzT+ujfmUKfP+Z
cdjsHN0vHOvobHhkawTMYdSfBVuoFP37+jEaFCeHZWiJLxGbFfrlblgQkTtDcRQmFAQOmAVp0mlw
GDju/hLS3qnyeJzAQhek4i/I+L5N7obS1pNQJE1stvZKcnlbh3aKPFgzvekj6u0l8JYGjAZ6p6Va
RNUNDS1rypKD0WPb8BYZ6PO9jkJH43uaYkhvHdTGFQJ9QwYCoc3v7pam23xgTN00IDnhPYWi62LS
sbhpDC3Pf4//ogTUWf7K40rOjoBPZuyePk2YrtTNtaIYEBPiv2BgIlquq7HUu5tGDDG6Hx+pWiXw
yVlbzYJc3HOq1NjwN68qmKG8gbzrR6kc4mmZNrUasDoE9o73OtAnk2TkB06v4DPpF2QvFrMTamyg
x5QBsJdm/58+2MDRVPV1qNAdlmNBxP4tgqqZDco+FuXUM04B74R7RmVeVnLkrPUidWI1Os+ppbMw
mrJnnUwt8TPdBJ4FoS9lOGafN+HSg9/CkjcgfNKqgk/uM/m6YPtZ3FeYTB6Ys1605A3CdoeJ843w
6+/RDKcyTJtZkPv45VaPTlJSwNJdA+4yZFYhDAM2fn/CWm31CKK6BgzjR3Ibf+YVfHtih/GhXvRi
9wRM/abqPQXxorHw1d+aw/rc+NFYPCFOgkZqFVT7zGCpYvhTAMG6rqJvpDT0qQhCK9JOTgbsoKHf
uNmtL4kCRX/TM60l0Gw2jI9ZJnS24AYKi+8ha/KyhlnawxdBPYV2hN4gWnzQHojQt2/SRx32vRXx
mYr9DyqGDzFQqVx7DaJPyVAeHGUV7103YckCVm9FICgmgHt1nx9ihGAcO7TGg4OiKYRH8xHcDbwC
3eFU/mOYNh7N6d0y+VbIZh7Llf5cTxdpj13DWvUV+JZmmhaWCl9ISTWCrpBxR51en+WzBHcq9jnz
6C9FiO8tHtDJ1NnFL9ZqaeEMiPOPajxATQS00lqXeGJ+aViWh1DYQsmKs4tK7IgzeA5hFVN2dIXc
A58pQb54/0cX0pPleOD6j5Vuq3w7V1vDDcvFuCbCUGuxi66Z+SnThrnTNXQ/fWrUdrBtHbRVGQWh
US/xfG3VG82INhlLroKK2RUL0ycL0ntsWz8RxAIsddqIGyLB6lcgF8gdRoMwCK/zjtsqjYwAFFmT
Pxsy8pRZrIYV7qTlQfHgCfLP9Kwe7rdRTDxb0TTXybIwVCAm3g+kroUr0WFvduxvpopAzOM9Fi44
LDd5O/ccCO4n+8NP8IVEmv1KNcMQWWfQQTdVz2SdmxAuL9jcy1O6KYItbxAj5/5lCl0Lw418mLQF
nR2sYu/9qNTeJj947GqKSssijC4ydVK1p3xtTdAPVCqulnbpp078UIyO0LagaGwxolWZNSFF184w
RQWc318tmKcDWyckZAbkNnaa80xOdxGYgnSna3dV321qnKpjj90QfErOREOPgsMYzG7Y3XK4Be/U
HA/0nhk1+BaeYAWQSCT40u6vWcvANJlMp9+1TslPYY15kamFZJFI3DFhRqM7AwJywSez68irVf3i
t7gBYbIYQMMyUsTRCTRxKc1tnrmcibC6EQSQkFYervWe+TB3eTQvvHk+vvp9gBiL7UiV2VdqFhZ7
GiN56GAiacXoS3lDN3KL9PrYnnTn78r9DysCDbYsAe/0So+1Z9+/C0waNBqv2aqp9jrPdRuezRd+
r9TqDWQKv49ti0CMqS4f22LK0rJjCAcZLz4GGyXrRrN1EVkwtUCMj7fJ3ItT9/TSMPCnPStlvW3/
FXvQhqSCJMiu4z1kHvSVB1zz0iKUbCq2783GPtG08eaEzGU/J37lS4cfXbyEpZ3LDFrzgPmsStP+
LZL+83hRoA/O3emJOeRejSStYwzzr7C2E2YzprjLDrR1lUMOviAlL9K3P1T9Q9oxgu+0wgS5buBM
fnmvFAutmQU35+EKGTyoaVhuqPZsckjJcyh8xZExJ59L018TLTW0xu3yyZlCX0Ld5gTg8fJyx2CE
g3rg7a0Ttk0/SAFZC7myZB3V/jhtdRVitwSLjBJHeSjzBQlcHq36uy8BWyHmOCOKE31JSWSit96M
azD6F3yajjTAPmKCRMOZGY0NMvSUw9hcUb4xHSFJed7MI74JPcbp2gauMbkAVRRy5PsNe4sAxmYx
qz9YsSvbaKH10z2fHGsN4J/b5LUFIaCUHoG7u+EQ9iRYcxW5wZnkQ1UigtsecuSW25AiIdNRmCAi
ik7shEB5L/oZk15wzaUf84GlRWKIzJcPyh11SA00lH+Wzcj+G2E8kmQjDvhbha2piCyfcoYQB6h5
m4OUnaZq3VJjmqUeL+/N5LxhjeOv1FcMwWPynNnbddhDPtsgCTk/d3V1w1B1zh7vjc9qFvbZL7Rn
BzWyykC7TM14kYZxkphquXBQnx5ImtFHgmm6OmOxc5YVjOz44LRp/B9NQMlqzRkMXf1iXJmhquuz
tseF+wFl8Fm7tTPu0e1Oo13yXUcR4Yd7zZz2gBjDDn5UqEe7XTdt8yEn9URGNb8jXDXxbXCd1bgW
2uTYrtLWp82BIdeaHETask1CVAks5TsTAHEgkXFh/6sYgWN7/wIXFwX6R3mEVUv12p6tQkItD/bj
E6G8sBP/ybqUnZP6W1V3OmZ4DHJelN0eQf2Pp2Nm2v3UrbFp1iKjhdrxuI+fsmuQ4I7vHyQmaDLG
caLjZZl3aSVlSq3OWxp+z2aLTFZgihZuFwiuDMds5a067CVMNXB4OzKFp6HZnd/ShdIJLVylefyS
x74045RbtkZhzWRYrROyvrdJ2UEMD4YYCQU54VN3ktAD72oKUt775UWZ5ACycvOfOq/OdspLs1Na
lOb7KOcxKTZs9Cq4vZCwFvGe7UStoDWcifuT/6cdufpufVWog0RqSrIIVJCoioCcW+fOLyxLYrEM
IauKWZ9o38vLfaXlKRPdTdWGUDbHNUY9J3DpsZSRuP1MABly0c4rgAEf1sKz5t8RFz1M/CVGyVg8
suWylYa0kUDT/FzuSpTjV0YR0GU5E06E9bkGpJxi3RaxV5DjJfGyew/ro4KcIHB7Hugtz7tzVlEs
8ViIURu5rQy2/NkgmPeNDlKUHU1yJWQnN+JDFkv8jZmH0joOPv7wOFoledJ+1ByXsvasff03p8rI
fx8liJViegdjKHukkJNnrSoe2S0H9u5oHtkMGFr+twLTu1142c2WmxEup/LwPoyYBJoUK762ZRaA
qQhiqxtVQHDCie7Oa0osp050pYvRXefkCvFM7GsqvHGsv8nFmEc59loxnOOIKncvZRQ5dueWyKdN
JkHmkYmKzc3pUaLC6QZqzoxLJb6XdLvGnxrFILXCkV/5LCvom6pKQPe65mRxyr2VH0e2CRlL33Bf
ayfm6955PJ2UzB0TmlLCqm5wh57FGBfKgq5scdlxL0FKmJ9n2va3i70yJx4wTjH6dAIXbMPI1KqY
c7GifpBSuN+HMC4t2PGyNsEMrQFJ5vGF7CCh9yHChx9dNkpI77ZPzvHaPsWuTjndocAKKFc/yqRx
VMY+idXpR1ORYWyoJZHQuv+kntBWsibAL/n0+dKZpo0ptCbMRu2a1WL3yvp1VSwRJUiptJgrYzm9
fcgPv5Dl+XMfxyalr0wbnHy/zEOXzd1wVQ6II0P6/NTZBObF6L2Eugi4actBFjCSfygbiR/erZFW
jDIpkpUm3Ns5sC3qzVlUuOBHJ0IeHOlfgg89Lcrah0WQMvKQEirZ1s1m/c5eG/l9f2y9deHM1de/
5z31ab+lW4myEQbE2Z65pNHnva2yn3xWXk+zsV4PWpjUCbhVfFo5jEAeoGMvL7q7H/A7Y4+okHmh
fUoyQilj5S9yxd2YIvOeXHI4piTg9XFlzoBSaAWfyMBd7D32V8voFIQ55G1R8nKrCglu5lMS7IPH
YAaMjZUh9fPfi0Xl4S5GEM5rx8HlJhXQYRdtaudLEx0evvmQucb3D0nj26iwW2d55K8JiabzxP7o
42KsiB5MNP3Ypstaohs368Xmwl3RyujBDSfZAke4mAzvYXjTY6M42coIuuz7RWf3ot6O4Q7FlNmD
mlB1vkuSieVxoCfT6BGdCjxKESJjQBRKgqpa80SbSZm9KAffMCouNeUIPKudwDCQAXBoTjJFkAiT
Gwc/q2w/BorCPAEsDLS7tEYl+CrfkhD8mggltH2sBn3PTZxLqlgw3Xk+t/vrhTlrsC2rFcKjOKkg
xi3gxAshm1ayYura1/m3f3NLFLfyrVSbTzFzajKNVjAsAQ0yVf8EBqrGn1qTLDKbJLAkAQpQwsdy
V7FblLb1Kwsuhh2TB8fClehSZcCINZVIHtcggTj9RrT6IclTgB7hga3RCkqEhC4I4+Ca6ZPvIAle
O95LgGU/GdzOutO4DukF7EakRQcZxBkfPpKeO1JAYIwnsqDWTR++Og3YNMJZf59Db/5/awiuL9XH
f7v+mrr5VFQxDN9oakHGhjhilkzsxjXfbmJ8vzxPvZb4PjjDaPdS7efCge+y1ntFBF/M2RMP93cz
Hc6OOp5Ah68UX+Uze6pmZuxo2xdBPcMrZA5O2/Qk+v8+IeMhmbdzwI5aud7QwmKxBBG66691zWqs
Ihx1HX35IsWV4Xt6Tk1GXCYGMkbD4mYGNafPthA5IBsAqqQ8hLK/J34iIpFzW868/8WNl2pYcpp5
sBKSkrC0FAUpYA/7PBLXa6ZVyrwmqNpV4WKFkFk95nguK8UZBO0W3u4ApbmLYIssp6Nk6zWFFV+y
xo+2mcuCare07mUj1KbZrQNe/E3yyzNWVOiadSfnBqs7mWtlzJLrATHldyw6WCRiiY3v7tVq34Aa
k/fQuwHRou5a4gTfmYTyFBhj2t8U9LutImeILRdSpk+UyQKkdAuhpzLSIQo7HdaOQMfr34D52iiV
QN0A19VzgX47RjBTUTGAUKHjD8CzGULg0UZRJHL4k079hKo9cUDwukO+dOi5w69prn623TJq+Sw7
TV7OsCZ1UYW4TwWYcx/Rlj5SaljKGC95Wat/x1LGzr17sf47JWmC9U8alZWa+QjKq9a50WIY8gmO
8N5biMKr6hAU8wVtLJK2YDA55mu7mhALW6gqq7rdhsBUPHBHiK6taE460RStK78fjJyP5ZSF0TkN
CTSXJs/lpZ7F6BqJGwceFIY5UT3LCww/R9szZPZYtbm2oUv76LsJfT0zJCbkQD1cGt6AVYx1CoJ5
m5040TBzsBqCHe8AGecmigabtZUX8z7yaN6XkI68tfITiOfwm4un/qchYhM9dlJoyqG1922SiNnQ
+QBSSqpsO0xmb+YIkopng1lLXVb2RE22PyPLIHoOcooGGTbUv5t5X8WW1Zutyh25SWPW6YL1W9ed
HjOaC9dJC+Hk04FxZmSJMnREjp7KlNMtksrW/s2290qDabsKUCsXrA+i4EicGy3HRSGirVA4HXEr
47M8KX/KX59r4j/9dA8NYAdDkLQRZPc3bB9xK2gUnkSvMKIeKoGT3C1JBQ11mFBTYbY9rTV9IGXA
8fMQiUw1r9SjMGM0VKOmDGr9V4vE7VqjfWRZN45MzaxIEEHhiJyOc2iHdD5CnAuXG0qBNKFgaKA9
w95YcHfoRixMq0BzzTeW1IwfzKjB1uCATQhYHwv5jtCi8nj8T9t7trDMZn/Rap7JIQSyWJ4tJime
b/Gh9iVNervjCDMHOtkqZJ4h3TXVfA1Lg/8GmbUqqpOtGlOi1DmWR+zuSPzK0ADhXdT7/4i3B9ef
r8pZNIcsDgG4gHNtNefo5OkI8+CUb7uWZrslZMSuiPSy9Ca1dzL4a89Cq7INHqTw+J8bLoeK+R5W
4YPyjDWsFedL/DbAPo2g6axKssELrlW/LSRZM1Zd4JmKNGsMt6zsrOl9GBm5f3soJP6lAqMLmVLK
2WrFJzRMQtEhCAuEbxM0nwvxCJjn2Zjfv1IetWEd8N9rfmavPCLNBfP67cWrgvoSJEqgJ/Ua2oxc
Pi36YmmMDPXGFdMGuySFjwiT65kOcqEVFhAijIQpyxVxMUEYT5A/fOb/mYJ8LVxNQptqvwUc6TQV
oLCxYXdap1jvldNWkIT8UEv+kMVnAwK3coXnGlpx88+fNWa+F7AgRQJUNGSb2xmrlkinENLAlVl5
02Fj9E9YD4iip3lPWW0gSjJjeuCtGzForcVfoPizvcng891uOg9hPfzOT1xwlkMbFWvq+HT8OVl2
Qvqhdq9Z5NBfiiIAe62LgsjUnBPsn0CdQsrvAud1jjnIWUHa63tpMPlb9+jQq1FOfnFs6iNVEmiL
tHM7F7RqvsAFlR5FZltRsAKh43J2FuWlN4Q2tPegsVRjIyTocby/bi3FCgQXIatxdguNJboccCGw
n51HP7ql9GZk9IaFy5PebfJLIbXp6q0QkX4RRhMi76u2aur1Lyit+JHqqUH4ORUZW71uKbyasKKe
WecKvLCQKDRHsoVaoJaf97CIJxtcuXEMFT7vTPMYG0aFb/o3JJmsRCeHJcihEwS5loxXWlaCNORJ
4EVnLSlMwvEidzkYJ1pzykqH7ha31F+203/OXgcFwIUzkfaAJ6aehsT7j2pYmZvoucTq9YnOFTDg
Zp0ukPV2kMthhwXFcRjcjgN3jdLgaaphVRNyFfoDN8kHRNkCMkeeM4712gNOktGkr1yTTjm0jSaw
RUZ2cab1qNq9iRgt4gLdvfmb2UKnDl4Y9kpeQh84dEs+T6/D1DK5VnLWJDe6xzhYh8zVPK1m42Rv
GELgta0WdcMkQlNLbCP4RN2juA5yhdNSzjxg0iPFV+jQzVXucgSWdUeliV9jJy6SRCHNTg6Gpmpj
0X+mQ719RI9En2l40K7EpWg/Dfw5REliJBpm2GAXNk0QTygM2Lhg11fhomFXb7zpWUYC0KGSLbJk
QD1epbu2NAravuBCgdyTdOdsCNSdgE081K8C5U04PmbB/13TvEAPE+5sjPK3hlY7iEi3YOgLpjzp
ZYs6nyvNPXHyE7gy9jTjG4L6Wd7ZkOaGEkITky+Es8P3CxXp8cRbePqVdUTNyL9fc9hQCgf0E5Ho
uVZql49/Lpd/Rc+etMS4eBImTmxVzQdoQZ+3ROohacjH/3Kh0DT2nD6ub6jsXh07B6+imhKU128Z
Kvodi6Ejx4uYK34b6r87XWNJzRRt31KmrHsUMicf7kwuIEz5+evgksRRQcQhE7uVzZXW4wjjxp69
9PBtuEOfmOzAI+knr0ai21RwrLHfugz3vTZIlUG978O9nRdaUwARlCsWa2P+aDZ2KExo5J0mE2AF
V9ozcnkNXppeZTkhBaqSjT+Fyb0N2xyT7m3NfxAjVF3cOVP2SXD9PRhQtav6EwCOxx3Gg3bt3Zkk
2MLiIt9/95QTcarqN5NkclCLdSqh6+XL/DDRALHRNuaDQMAulZq1VzmX8Fyb9tFY+W+9+LOc1UCU
q/LTURqfnq24RGpDgiLBLRDVlicTewNoP3vinaO/gV69AZ5TZcq40h0v1eJfHg6W3890FrOR/Iys
iiJhRfXIJiT/H5rIK21x5arUja7OBI5yJMH+mcJ6b6gUcsn9hqjX/X1pvE/r3hewD+1q6o+E0qXC
1995W79+MXcibJRHIVm2PjHFGy1WCai/mjhx8yi0JQaX9TE6q9iM3imlxzVAWIpg2bgfnfSIxklZ
+/sk/LMqIl54DyDvrz5w57GGLKzBasf16A/IprVmeas8HVgJMtqvoW1MwTb7XWd1B6U5LsSNIVNr
PZKDnYNDEnxXNQjyz2hYF0ljAWgXyPv4UCnvx2ycuXJaeh84c1qPKOHPncVDxezJHfdNySj07FUm
gvX17Lq2XnzgbJkbNDnehFJS5p/YRZB7tIsfi9wxzYNzPG37PKnsJ8I9O5gcCinoNYoA17VB+hIz
TjmmTIJw/zwnNr/enKyrjLb8wraN0MLhcrUU3Y/BjTn6E3ZWQ3SX/6W3W49EXT69Ik/n8eRzF9r4
XBBF9Gf8S1Gu4pd3ZAfMiOcxzfYpembusiDVmXsFo5bwnwvPOJKiGWnimNxMZ1J52BKQKFSvCkYu
8/LnHpIs4gB6eBp30ZA2b0HuQqfyY4cH49mS4l+6Yx+iPV9YP46WAPHLG+VJnXrlwAHohuiOnVN3
NAEhunZBWHJpzHyBgesDQvYoPNXqbul1ART0YzvAp7TpcrZKGaT3qbQz9YGtomvAakyjLSs/t89x
WxPxrd2pLYgSG26uuDLI0V75aP2UgNlnaHSNtrMiSacY9Yf6W13sro4Bbnl8UBRa/EbR9qM5Ml3I
tfYC6ivMt8x2TKCk1XVYJUMlixTiGJDGHT6Xl+s9/6E2KO3tFnG8ySTfPJyETxwb74vlnbm+vnDP
uDcEx+c+7HyHAA8XnBO+SajmcbJjBqRFJJe1fwv04NI2fVjezYyA/UCceCKS7MeXXLeO5aF/B0Zz
or0Rr+gZhwCK6LhreUvV2hHiHZFsPYamW+Qb3avCdD67YFWziasquHtJGvQUV136dNdXuWDr8UL9
Lgv3DzMXXkbDit2fAbD3lKmwJkhgN2iEPJs7FMi8InhY2p+sHqGKomvDxGZb2YFpwj8/10vqYa+T
w3nFM70+O7wScnpzZx8eedbmte5M+JBYULE45yu0FCmAuqoGaZ96FbpqBS3UmAqi4+Y9Dk6U/Q45
oebhlizHr206O5qKtDU8w9Ej9RpeLV7mmJ4++EgxlghS+KCiwGRaSTDnrKhgbKOivtE+AMyqnCoS
TpNw1JeAPdTt2C4sd22KPrsRhncyYPCKkcDIyAXIbyjf8uBupAmtVylXn2MREtc+cm1d4cgwhE6j
xM583tfp6fzjwr1zsxR/tiqnuW8iMy46c8+Wb5/JBd7pEw/wTKBz9U2IT42etLn4a+9SycUDxD3s
TvCisAL91MGwK++pHBE3C8H1nle0CZKRIFNDOy1iD/4ynoZRDEVtamD5PDlAywddhMHulRRSYInl
RMWan32SjVTI+lZW9AKSatsp7D9Fb+EGqrob78n7CVBve3BFp9Id8aSqniGBJQ3Nk3KRY1bRyXh0
W0J4EqWRl8rUO2tBYNcQdlTYiwwiEYe5Zu4niwysYEkgEvApTcIhX0LL4HOyISIqa+rdysCLP1Nn
vlinncgVbWHAZQ6frgWbQap24wfzpIgD/2KGnHvjNkP9APVpF9JfoXA07cbQ5GwKagaUkdmg55lj
lEkIks9yZp1QBvReDoAr4kfaEpwfYliIT9t1BRyH0nju3YYQxt/GtJM+RotH/UtY+sBv72/6aFer
WcUdZnpA2CTODuuvaBxY8xFfHIbexS5YFuTO5du07tFUy++eB4CL4N8hQ5m80AssFTPc6EE6WLjJ
F/IVFhN/b/I+FnzTwHrv86g7KE5D7sGX6yw7HMrSVXKDVVwFVMo9+49H2DaYVtCFTJSyIsxB+9sN
kE52kYU+IJuYcSd/MhmN6Vlix0MXqiShvOpiG//dLVL/F/lvfK4y4ooypFeon/KbeD89h0pYQP1f
Oqqoz+Gl/k1QKurtFuQYCsMGAQIKzXg3FENJ/+fdqtwXDdB+AQD9mWsS2LDpUGc6QbvD3svTQtMt
GfzD/Lf56Ncc+Ty/7qLxzHwGuVYHnjPHGEVBoVC/skiLsslRRuB60qfJa4tdhhuR+D62THe6WPLS
93uTBzox3Aa7hhRblDwoFw7NLuvOOKlF3RD2xprDhqyYV0I4BgSoPwPpoW+to7+GBUuDMKx0Ftpl
ejlo9ZgTlvT77a22XbocqXysPm4E0Wj2496nN8h3TjdXCnLM8SvYkFvCTyEliWs0JZAmrvwtOpty
x75AYiIH8ZS0PyXW5KRkjTasN8BEHWvTqOaiZKloTAlBwNmw2qfCUZx6/65vukKQZZKV/9i3+Cra
+xZ+ZwvFmhL+KT97usShXIIigDejsaMyl7aMlLdJbB+lG91DoMPFQOsw4aADnF1JncVNi/UYbaSu
NAfXSmJdPpR42y6IkAvAIWizz2XzbIFP6LRy8X2ZHhQ1vdrMwnLFEBJKWvZfUspjkBLgKDpWQKpQ
AXq6WwKX8U+BEp9BYUUwc056/5Y53WxdYbK2lNHDlPIXpkO9E+vL6Y/zEAXQu45fdo92HT1qQ90P
y97B368ySPXcd5kFqESTJtWjyFwkW9H60+g//wjxAJcZ5FEUl0uUGaNS1xjBD5GIejcWJbXEO5nZ
uRgLi8VH7UqL83dwY3z9ZPzU/EdelBzeZArXO585VmAZQAHtf1xBKBiKV/42qssSr6Xp6ORAiYbZ
f3VhvnGGyYtkMtZ3vA9QKbqeYNhjncnCypx0x9mW3hyXtHNXiwgTYeHwcXCJnFFEuP0uwR5FvXjh
GakT2rv593/vRk0SbCrMHeL8USyZ2uHTTKawNaRNjGVVuupWgayE18tUSX9UBaT+Ug4I45SMfwxn
wHK8L1oR7I3oGsWSymQHkDP/Kx3tQlIg7Pzl0tHwU+1RDIogpW3ABMAvVtFJjSuAAA6qPhHaZHKA
CRUge9sGK5KSRNxqTeiJHQ2FYMYLgCLy5QZxK4l4lWPyK+nvmr6EG1BYF6Lu21USrqbnkPqqSoNp
jzBaUowxeb4FPhovj91yc4dc7sNkcpaSZySUrztwt1P19XsVz0iE/Lltp6wWbHK76y4teB2o6XgM
qdhCfCvy3h4VssKVMc53coUKBJbnAN/udcmYv0aqc5P4IiCE8Bsyb0kYtsl6YhcZ3TH/3PDNCiP6
9yk1alwtXXHaLFJnOjhb8VmZ7xtbbnOW+Tc/LK0RUjoNA49rdaf8lE00MNtqAjnXQu0YmNVOpB7n
D/Ri6uRQDXzhpmU1BX2izPF8ToclukJn6VSJIYylrc9xD6w07z6Rcnsc9AqtBuUpRCfgTTjb02Mx
W1KxhqmbNIMpESdANhTdFgoZpJclQc9QZx66itJ6e428PCK3maorbb+h/9kihpA740+CXe2EYnIs
t9D/TbGWh/PdHD/lIG7bTgYFDJ6o0tnrroBbPdKehpF6ZL9+Mr6KhZ4zKqqgzmtakU7TdSFMVmeP
BDTFP75KvEifDNDxcub1eF6XnA8tkihyhVd42Z2vDCRLcm6kiuVJDqV1Q458Q4Wv5jOlHLAPyked
pCC8iniNYDwkC9XImXHrJNPYtkgYE06OVL5exCBknQ2vUXOK0BAsfXBagiHQktoqpImdJ/Sww/AP
3KQAuTqDeWlkAaG129k8hHEPOt0aPpxSTj5rFikqRiBFcBAKPuneXcznweS7ok97vcIhm8oDpPQv
M09LnQlCX9QukAioz9brAlvi27QzDsDUGIWCJ36cgQNCjyFzKr2lTKRrb3Z3fLUNVPXcGyp2YriT
Y4Ce/6/I9FNJ64nLclLi3QW9txrdOZxwZnlKog2nQMAAQsjiK5za+H2170HWb7LHP1IXHkahYw7k
qzMnP5qTd5RnWtbjvlsTsJ6ffGISeQjV7Yo0y35wFImVLj4crbO4N0tfxWemax0HitcUmaXlfPcy
7vK4i0eo7z8VspY6ORbmSvHULLCluQDnDDlHT5Hk5krxC3uPmyqNVD4uo9RdokmRgGM1atGhxgzi
cPMa2pb9dMeZnTKQ49jGToVjbvHWJr4VhYe21qLrc0bbulDePfj4bw9c8YrYFeBgEfCyOBV82HJ4
v9/XOCRioFOyW0LT9Cp2l0JuCAzSlS4TxSWQvxxtmI8JVfm4rZ224gjT86Pird/JALE7cHBkq26Y
8Iuwi6p0fEY4IwrOyzYSi16el+orniKzmdAK+VWd51SY6yShNma53JvH8KIowJgCIaydbeEhl2TT
QwjF+yKa3D1OriPzoNkyECM1xhfNstHY7f2dHWTpHhqVnWdZhN+Z5fJIlKvRu3WFcfhabDoNPmTV
y/bg3+AaSVqyOWDbQirVohQYy9+9zK80tsggehZgORTAFGb+6GzDiARWriNY+LkGMK4RpoTW6Srb
xiTlj1Ii8u0Ie4gvYfYQOef1GNw3Zd9wTzGXXjL2+rY/xKd/R6uqMhH+jGvTcB9ADYjEbYGdEC40
kYZs6diGrhugs5WQFRdFtOUMcEn5dq8WNIeyCzOkUhyloSzVCpwk+VKkWH1aGfwjZR8qYe9H3MDm
UGb8KeIGhNNB6yxnam1coFaHLjCE3MFrkNysaocGhHUrUXkaSOkZsmdOwOpD3wh75gem68/VQEWI
bBT+5FgoAl8yc2TGUGqUlK7xJXsM2TDK6B+4g4ofsoFUTq918IN57OM5Iqj7y1FfCSSH+UUr0pIh
I/Jgc4sl6LcLDtOwPyhz01kGPtz7h+VEnCydtEu2OMZ+ZIEh7EHXymGpYSQibY58BjGiOxWFvPu7
T8gyoCAXAX65URl3EsGi06DJdBsmBz1afI1YTx6zpvuFGnYPngpf0K8YE/7e0ejXh9WQ1f2iXzIK
PSrMkbIlS4D9Co+JNnp/xlBIHIrLh2LCQxqIlO4QWx57qwf0bmp8ltULhtQQ6CRdHYvB9HJdrPr8
wb2wyhCMxzP9NBfLpE912g62ld7m9PF7WRJi+U/un6kavDT5/1LrfKXIrUAXX3Tq4V85kB3vuGwQ
/ZRgdB88xpVIKct1l6cEuniUl2sI0Nn2Q/gUbA5TWcJJNX157SIbaucQj3iKCydaN0SKAzPURBj5
IZzDasy1LLT/nz1eeViKSyLnDohBp1pCPrf0elOxWG/DDtL2/ztqqmJYdH5imTVYchJRMKyLCtkL
Hm45Bj151JZnfMURYunTv3MsGnFiCxzhbP9EZnXoRSqLYV5zuuD8tkkfthL2VItHu/bLtfAOEgdx
u06c3+bWHY2EaqvQ7H7yBLja2qRa7ui6KIykMgARf6FCW2kEUyE9qFgKNMcqg6rQPqLbRmcV/xwc
jlcGtzpojn9VRsdKMXfGyhO6LSx1d1/4J8gzW2KQeNdHOwW77S7QlnXnv3iT63jmPn6nKuWHBw2C
44H1TsxqRpAUWDa/DOYLCGmWj8lW3vkhR0+JrtBoOOmu3n4twjkQCQv5pzaMqN5MFxeSDodERRNp
Q9gMtAFQ324gydFdh6/7GMoY6Aza7xPFmz0uBEorogOlJP2BNw0THEEWk5zIy/doLrkU1VPE9RN0
lYll9GjXZ3deQmWZVwC7AVB8hVz708pnmRYxExbDjgce64g9KriSsvFguXc+wQNUDW5l7HWDcMAY
JN00w98gLulyIdfvAFsbSgOa0tJ8DGk7WAJ7orx8Oep86vXHl3DTpvbpuu2vpnHtz7XADF1GxH0L
wDEE5ShHcFxKrDMN6CyG8/GXmfQ7trGib673nFMQ8gi8xL7K27+qnMQstHaTB0Nl/Pj3f7YMPeDP
2F4e4PVtuv1FxBcYCozFcVpjMAkMJvN3bJTZIxV7QNXO97wSaqgA9dSvlj3RsLmBleENUm0xDwEg
T5ZtHcB2LWsXMwIgSm+fs7bro7cGJoRgrFmTaR9Z9ZrCFU/YUBuSBjSEJF8HUYXTbStugAnJuWFh
6AcslUa+8GDE//oO0RPaQM+x35ZkZhcZdDv9Z9FTOWFll2NvMzvYaNjaZ57HygeB9X6cfAiLINN0
8hRrpEd69K9xB978ldAUs+el09lC5lxNJnNaY/BCDIsaouvSFL6eSGUyQzg2934PzGZcGjFCq1wp
pE5AhsO9WYiQIKrAbHp5HoDJOShYkSb7I8pOpmjtBDrUpEHn50JhS8aZH2jSlyCmCfx/OUAWf/gR
hIiU6puskP/FHXk0N0WyDMPtZFdqrLXGQR3cEeMzVea9xLmP9ucVVZiBf9MM2C9c2QlNS+vdeD83
rh0R1LF9aWYPUt8vWm8iF9BW0hZ2PtIGZX8VqofPBgetj4QmSgBfmh2pfyYmOOr5wrdlOnG3d23/
i3OPZXuAt1N5Mx4LYjSE+yd2AGrDaxXoj1zkjdcbnHCX7j01E86SG3CiJpYoJWz6pFDY/BhN/qQ+
ws9mNP1vhDoVuS6iXYjUmYKa1IFyhL1e19EJUb8tBlLn5QrqhradppayxQz2FJTptn74R0qmGc1j
OWGNeXhul+1F7j1D6Wia0jdSSd9xeexNbNYiqiiz+iHcpkiDQLHQoUl06C84tqfYsmqkA9XAJIBC
6K/AQjfo34orkSkSNHO9RwuehpMsSU0xWwTvXifQRN2SFsVm4/SkqzgjW8+DdSEmubuE8d18ivKn
5txc8hODPerOa0K8E98IDFVCYmD7T8sngYBhG46CHYiUbBXm+uBWUsxvGQ8vhnesL1l3Ua6Tvybl
uhxa5Zcuk5JmQPMw/8lC6BoF0fDz0n9nmOsttME8XbAkbCOSNtyxkuOcttjFWJEyLEjwA+OhBcTa
qakezgj2bREDdaTPB3mzqSJO/7/HYnHRJN5NVx/Y85jtLlf3i5IbLuMHz2Jw/FalhPuMjpld/s70
G+JCBKjQ0/yPu/Xl0sVeED3tNLQfH2wBlGFPOpK9ZBxP9K7FjNBCINz2AX104M/lAyCkci1T0ULM
6pd3GD/miwLuFlWqOi6EPlcdh2h7y7uTWfr9Y9jPqyDSutiHnEd1lTUuMkEk8miDsTmiLoah8ung
VJnf6Xp2ZyFQ1fEgEZPS6WQ29uJbujWZ5y272I5/QaMywV9FhDS/nR0wbJB71nin6mZgRS5xtLdt
Yzn6UyCTmitY3YNFHlQz7kFtf9wsCtnM5Rh/QvZaYck1seUrIlTrazLvFvNH0ASKsHY4wreWZOGA
OTxEfrsVP7xq0+INxqCM21ZoLInqbfmffwyocMp6TcqHqT/FvcjJXLVujx+kDBL3hAzG9b3Y0lFr
O2j9qTFsa4b50SKfzhPIXeJr6SwqA4OdaK1a/QgTwici3kzRpzH4pry2lbfSOxDSviorCKgF8clB
uWhsf+MmF+tRetcGTFbwhksG7M5Eif7GtYxjqh9hUSCXgfuBBNQI6aKNb1whC10khNdl7q3GB6Bz
lwD2a5gDXUZ0kaExfs+02sEltkMtXU03+qNuHyZ0NUifk0GGYbNdPHRPatZUlzVhR+LR4G/6Ki//
Qb03Lxg/g4RFTebsjUsH221O0ZL1TH0+LwMQpPAnE6T6gNHC00l5thLKEP0+uMsEDBkJwayU6zCM
ZWkA+cIhM3MrYdE8WpNHYm7nDWPAAtP9AX6y5fDlIqLPZG+02xkGGULjV5r/ltoJwNDjHYqrh0kW
ShuxjlOD4R+GXjLNbA+UOY3Cc0o2feLGA0O8ue/yG4YzYl3pd56ELPh7F4i6klhuI+RYrYkgsRjw
9unZaQOyM+RVLAVk8tpUnh3cy2HgOHXRUPc5TRB75gyf8fys3fossvfJBq1vwY61v0pgQpK0ynHd
y7tWQYp9mvu8gX/4A3fJfozDyGaDyAERqtCF397T9lTgxjGhzxNkB2E8os4VdO08/HqwtFs33D7S
J6IuwzGsNS0OGuHx3jqwa+CHdq3hkc+uqk3Zek55EsUDJfjMbYZtN0+lgnB8DqEOBEQ6lcLwzcdm
bhJcvD2p/1b/CdYcZRLhpcD0XlvNazr21WzXK+gCrJ8sqW7My4u4UOkOilZz36MPj56Uf525DdSr
nJXvZQ9YN9VWG67htSrGpOb4Nwc4r5gnanUzI2VZMtCBbmlY3mZWR3MfZp9TPmvcd5kUaLahI2Gm
5Yz4CXW5hz8mTtZZwNE4H6Zox2OWhC22SCTuZwewpaHGa/zxmg6F97Ta3yVLKlgq1y7B553g3k1q
TITjIO//Y6RV8nmjwhBgslqQeuXYwaSzM8G2zHpGV/L1dayBWxtKz6cZF0fX9qhSUmVpdRqUx2up
xuqHyEVE3ucbZLi0i/LBDQowisg3p/mHeTFvZ/P8lJAvUDjF5I2af+4Sm/KLlOWhHiAPFmdHmfUw
i1axaZ878+yHCZ4WTOQKLrMUr0sq4FMGVv0InPGHWU5+jP4TUNrHgEosM/dKvtU23KlxQgP4mMGj
PnPq6oJsDVgHydEi6Ir5Wu+Tw9BsfsQNhXP7HC7DHVqVYNCXg1UK1h6fUvUjY5N+4ZSOIwSrCnr+
KIJYwJhmSHWJ1R6R8NDgGfNBCZcm3bcvpmdDfUd5H8nkTb41PbS2dqT+fyKQdInLghznI1Z719tX
ySUMrpiEQZF6TXR6EdA3rF//dy4neuRFY6wbqMMM9mUXo5JOsnML9OW3PooFQbKY3bxN86DUgIwP
/aEjOPUKjSQuxiSQov/bSAzppyOVIn69+eqz1oXNFtCxh3GCV+9RQ2mHE5lA1c85c0zoGr/Lstfw
efQ4HdIB1gQZEHSWBU6IqDznWpu1pwYqdEERK7cghZD5oQ2PjQsZBfiLlrEOzWSa03JaEyp9uQ8Z
/M/8vA0FMwU2SeuJkmYslls4GljuHOnHaJfZjtv6cg9xFacKeYpws2CFqKFwXAQSM2XXLlQkZjOh
R3Yn5m09JSYZWB419IQ9fjFMJu1+568P8c1hTrEmv6uOp6YKrZyQt5njZD+SodiAnncF8K21tQ0c
Esm3WyVQzGIalOzVDwv9/YF3Q7EQcsZVVKXS8uV83h4y+bvXHGKzXnYKp0To7v6ZGxzJi1x6fZyf
vDfIoArFuf/iPXAv5EI+76L09oX+cAXEq3tpQAIrSFLOEyTfVT6nZqWP6XD6e+d7r66LPFdPt2kC
4xwFYx2MYHCmhh4O8EerwtE6qOCeBDXqVKFUdBaY+2/QzVgU5nYJWmqzPnuYNCjXpLzuBE2vupXp
8N8tzLatgI7AGuD9y4xyHL0rJfiRmJSg1EKm57Kz0bGES5UhWugDd6/Spuv/eZdlgOqQ1EN1z7Ox
wxKBS7B+D1dMI9DWp4uihK4cHxXc7/unQ00jAnMzx1jZbk9Dm4WB8fti2vUDYAsrwSSYeuxEAoov
QzsvmW7UosLfvYjudLETNv0feWdwoMtm2itBoIbFY9GyLSUyvb0n7nGX8Fl+tud2jTmOc4fQGtGu
5FsoNVPikrylADpzzf8y1337cx7DI1N8M0y/OjLY/EgmPUPYtQnBVQ1hzJr3wCjk2kwxkvfBSnyG
xMlFEVi4gX3NzQ1PeQwSAZFY6Fjg0BINJ7NmrxYpyr8+tBczLGYYmwvFaTv+gcMZCegFU6RTly7Z
rS7FSRi3XFgliOX5gEPgxjvl4O4Tz2/+/Vcp21dw8WSOFg39QsOO2wKwZZyMGQEMbuVQrpd5608O
wesROI3EUEq6Mo2o9COueDNPOT9h+iCFSrU4SEbo2cnQhehYk+aij0WUDtb0UmUEAB0dOW1WVJ8h
orfo/1aawR5r1U0m1gfXJS72VmpSiW1YLlRjX+jhSxu4N/AOeGUCTaXbX4uagppOol/b3ljirG9B
f/Wou4K/7Is8REHfNpqyZXnc+BvNSRx6hw2944xEks22cgJIf3oRt7JSHG9sTHZbpBPXcqNeE07Y
34vMQEsoAmyo4pVia0D0iuwPR/filvNpNp1n0AhSunXoprOsn4Rt/W9TFVegMYUb2IYjcifMJUDG
aE/NDCvmvU9D3Y8mjLyeE5LN5bN7FGvCytWlXZhm+Q+Kjz4XLAHE6R7zFGu6NsY+upEqLL5CoVpj
8SZ4mJT2RV7vCtwErl2ipdKtfn46CuhvKB8NhJ1uOpDjhktNzKLFIaj/8AaMl7Le/h2RkxfbOCu/
+gPyttq+QdJyPdcxuDikzJU16tNNC42YsgjKHdVU/L1q8kJM+AVD5x2eTrnEHcgRoDtIY+2ieTkC
KNF28AD8p/5dRRwkCd10fkI2e9JXwz2mdk3KdUrLM4MKANrBwW6h9XOxPQBdJ+zCkJefh+Chw3h0
DbIJECBR+6e+lCXRrxgHbAjgZPJFm7jEEVCeUE4w13TIeJ+2NgSFaXukzA6vQO0vxgJi5ODoQRda
MnZIREgHYZGLsY5rexZwG2kUCXql9ilvtQ9YI048kUfJCakSqKK3ZkYuIMQpVVPyouRnWBhkjLyX
chsEi9TPQ8BfpqFNfOiHWfxPTMS8Ctw+qHmWZCCmAq+5nDUTLmBHbq7hbBBJfy8RKgrN04uhcnIH
t/ads88ByKiDs84is/uyU3GCq5dqhDpDBX/4vZaOKN0GnDAzCzOO9tsJEb4Db/MdBxg0Sb5DyraJ
5qxa9AF60r0LuD41ctbsJl51CgizdkwbltuvLw7E+FpmdNFtSxhLR0sHJXY/OdUnO9FzXmMHtCXn
axT1mmeY1P0d0BY4AM3nwn+4rv68LPLHi0REqUPjHmswJXo07vXV5JLRDAa99V22YoEOfzyx591f
nOZA3LLn7pKRWtVvb/OjoqG4BI4zPtiAz4kczX6fxFLbXg+d1aicf+WLqMSiK+J90uK6s7dGa8lu
Tic3MA6sFjCrtQYltV31xQdX6RoYcF0Y+urwWOs60sMLiqfYp7/z9xlrPkODg401OMsuva2WUaNv
H6BpOspnu1Px/3EbxO69C+L6iLICoS4xfTgTBaJkfjXupPJxaBjE2uvGPVRP8+F9+4GaxELtHdNC
Uy2wdsEMlTXPULd+fJUnPXXmB6vzP/rcQUVR785goJRUA7F/xAy63BEFDNPaJmvocIOtNSJ6NgpB
mPApwnYuyjXcSqzkPGZnio8skzHP9bgWf2Y18SBYm/5vucth9x4fCSTRpMPmxBjPweym6zcgET9F
zT11gOHm27oz6JZWzpkhAC27rURrI4MDkyNU9ZQXyqS+0cDGTp85eZOps6aluL7xXdYYzhHd1ij8
89InWX2s3Nk74lSxXNNjhyg4Xm/EYt0DKXMssSJjVUKjQA3DeJb73SQcFYyXYr+p3Sg06Ls1fViI
lxJJElYT8nVSmO8+/wSrWQF5Y68H9QT36ptXUfSodnbvLF1ytjmwtp5bMlMr6iHIn+e0P+p5K4Lc
N+khx32D0tj8Znjtl0HQor/eJ/pLdiFVAJI0wwPexfSQZ+3oNTygMjMW58BLNR9TP1L1a0REZhyJ
35ypnTDwy0vJjvI1DlNciW7Sz6QcBQyESPs8TWLrRyja13YvW3pvoJCEYP38TJEz0JvxInYRH/WK
vJGmZk4xTNLY4NHNzM1rgwQg0eylSo18nqK667cV+ZMng2cbM51hHV9WWC5/cffkMrD6Wpel8I7Q
oFTYyq8NY0v5xk2Nm+anp7eZb0jR/QcSWSWbnt/NpQciqjP8DgvSBQzpzYBySGWRwRXIvMk6pckt
jztU7nUbv5aCQ79zdKgWviJDmjbzziw+WHz8ysqaPGnecF/4h3owGiX6xkcZyo7cs8kfRDQEPKhD
ABz+o36ylv977LHVHI5qww8kQ0fRKTHYx3zzcBiQ9yPbGxyDvsmCSzilTAWRjyL1yRc3u2x2qbIr
MUqjfI3txaqnMwAMvKrKQYek523G2SxcghmBnrPdoIt3bky4CTu1zkcZEP3jSX+J+USiXJfH8J89
jzOP7tMVM0mAIbw5A3dBIoJqRZbL3YamRo1o82LP0NfQ1wEWqG0BoQO8b8ej3FYM90dK5HELLMkj
dOzoLT+rgO8MPromiBEIMl8+fAQgImdi2jTxJHhxANBs3nIR1JnyP/i/ZvMkgRsjPx4wH5zKueD4
quwyWOwRlP22hZQdqI6luyQIbyzuyiXt2QFWDidZWN/GwM+OOLpT5ITCI5oK+xB9jDOhb+rM8yT+
Y8o/Gmg5QQ704Kf+jZkfFqLL++c7s6uVRk7QA8F+J439IQCWe0ZqmGT+tKCFlaKpRNH1rOBHe8qE
yFyEpSSUy65WLzn2io6rACQwp7ujHpTe/ztAC3+Yw9E3BRGF2KzID5tPzhttwQdtugdJDNlz0Bx3
FLpq3Vx2pzJi2UpZO1n0Pu3h3Rh/nZLEg34MQw+267EqOBRoP5vBziBekho+OsFsR635urwp24E2
3uW1MJlAlHGCZ0RgAnapTGE1mfsRUcmDZT/XR/D0KS3zuvD22b3qR8Aq612tT9PQ7L0/G/nlacDV
/QATQ7FWPkwUeI3ei9YUZtL/eMj3+1ZPOz+LUGLrdqKtJ6J0wKdByeowWbx+OdECvKWVWLCFo51O
kCiOdqhgc4zKdLhSIiA50gxuDMKpQs3bMl33jq/jrVZuwavOMA7gA1xiHwq8APWfWGcEm6fVKF9f
oxt8ov9+9qJfNAAp21EYG2LVExun4R7wY8DAf4SvCVw20JVZdLNcX0ogBr8YG+Cpie2ncjbK8kq4
/zKYJFgCEpsWUYvFfe1xJ64/eZMTPR1U7WCbhaCObqjUZtLXMCNEaGeijkdrLlqilkukMmWY0jce
JWj/ozZWB+djJAj8BTv3PQW//IGeHvlvGSk4LOnd3vSnpnWeQlyA+zoSSazPUZX/8qETQQDzs07E
chage8pjpn0U1PcMlIkTj9rU/6AG1/ACkONdCIdHr+xL1llWa7X2eLALR0F0viP+4S7r9sQcKTiT
bKZ+xkGpStzb1W5WxBLet+9rMwRY6Yf3C8hLeaX2J+M9/4TY8xQQ4YjFdgpPCqLsCRQJA8Qsooz3
4FgOCPazS893YTZBH8IMGRMUSKCtulYgOLhLmvsvd0J2IC6XqkCHx/HJyPW5q5biKfAxdVECJNgw
4TSzAQSDyKFsf6QZ13cCpVOv90mrAlmEYhxSrqWIAL14spUGLNNPR/q6GwONq8Tm5OqqB9obvu3A
ePvzqMHfe8niBAB9iVs3Fyz+jPq/KrN1OWUUm6zodLxhpbU3NqRbCu2nQe2eG9iG3D7fT6N+tiwA
odIVMtQWYtkWq1icLodITyrPgDS5QqwmwgahzeeFyONkYADHFBL0eumFxmMdEhQb8xhXs6vEz+3O
nlHGRJngUFOtudSBRGONWh40Q4QXJJgYY3RU3KjzzYG1aa4s+BivItXKxif8zIe2AASSPMDoZwhJ
Pq3I7r/p/aFpfSu/8cR8BvVmYn9+CHDHYlv16L7pSUhbW0P3mzjd1dnD3mkI2ZG3isrRK+qITk3L
ER0tnU8m1YMBgPsXhXS+snTHf/jNbgvMSEIok2PgOW3wLPgTHmCJA5X0yPbdCvsEDAqElCM9I6OG
cv50M+t162qHzXUffG6ThYzGcvDPyuUONqCCBjm2WxIXunDhpTvy+Zf+XsHWBL2p+XJFzhpCmihD
i/iUSZv6JKfhNeOkWpmR74QEI/bLecIRPS3GmRAZZiRsZeUhirjqIBAZ6UpxZMu9TlQCWDwW5P/N
lsefnquitUf9SBLa52ZW2syJBXCwztKLe1+I55hemfDA8qpc+EN581cufJI2KQauif9zqfzfhVGm
q3yBplCy/cdKBzPqnEF+GiAudPjhuVhuMuIsakuinnqKDx2g5qsBxhcNjtQRDuc91TgCrBQQD2QF
NLjTD0Q4PO3Q22tMzfGoeNIIEk53B1kr9xI59fIH31wrwKx49eTe1YddbyR+0FLBRI78cEqLyRbG
KKK0J7AaNoUH4izPPBpy6jW2jBujM8zQ131NORbJalhwN9Cd5ankX4+7JhzW9g1Ry4C/XZXd/iom
TjP831ulVqP1qpFRzqIuJJHidBq6Rc+i0pQf4sUmXRJ4WM5UZiPGvR4Y2eT616GAegxKbtmaMbe2
CFnUMGi9J3ZS75c73vJXAkzihfcFJTatS9WhAoxVngdlOXkcqqUBscobJ5GyuekOD5AaUHTQ3QVt
hf3sN0vQskb1I+ShligT0rXV8+HDYPXdaRZBOPBLfMigJOMuw0X+WZX6RaVNXC2ZHf9KzPe23DXY
5LfJ4lTxNv9ZCK2qdjLbkiubhd9dUX/ZtC9STgaGA18AMf/odUjHHtYLsUAPknPTfSEGOTbrsm1a
+sQe77MvohwUsAn1BSrZzv3vS5XyXmrXOcqTAWgGlSvDgHM9v7X6KC8UgSTIHNqU+FPvdDoQwWlv
ua/Aai43vCv9tQ4BCPl0xXA4hcNAJktRM8VptHP4A+Wz3HhFb4brqKCBnCPBkQpGHUrkd0J6Ruu3
HDA4GXfoNZWJwpSkV4o2EZ78Jbs/5smnp/WGxyr4yqcs8z63hpgicN9h3PLlUqgGC/q7+0z88nab
fPHtwGAL2Fl/42Rsi1S9NY/qmySU5bNzF52r51uJVcKCrPxs6BX7YLXqYmscN5NOIQvBqm6+2Cx2
4DMfr+hUKvqAEt+nLtJh7xqr5hCz5szUKya9dVOLaEFn4OnK1g/XrGcFX4Je8G7kD3T0k1qqByGZ
x88ORKm+pDQSSFv9CmqfbCAlSC2dZkox7P+a/AucCi++pVuiYplE+ryyZNRtLzyPe5jsQQLr7k+T
1djDm2JC0GM6JlGVcTD84pc8hOJFmiXQyptw/Jsh0rrHhYo/bdDPtyL2+LXH6CcyKFWAgVJAco78
1NCYikMnOTgUS2t0e7aUk1Nbwk+yOyVdFnSdbe0VEWnw5fGhJasBzo1dOhLGGoken58R1LsNLsgp
NTj3sxTKgaBTM90KkBJ/8cyoZnKTMq6G7ohT556L9zaQYm8iBVoeNoQp0LQ8JCV6gcdJxdvL9JOu
JrVsrakONsS+FMa9eRBW1j3lmcrP7C5NXw1G0VmCq3XOqccJLHuIIVHvswtZQP/onuS2gkdvgSVF
FRc3fMputsSmoOUjctfgA++TwM3rva9OZpTrvaRzV+arDE9Iv/8DxcKVC0M1XNQpALgBB/kvGZRc
gf8KawrkV/V/4mxfD7ZKTa5gMG/F1NW9S9gVu4GzplSWver7tqrWlOSyFY/K3gAqqC1CBvxKoGRm
ExlafFKS7dEyGzMFl2NYdzV+Fk22r4IuObYSpzQahpJmz5x3Q1Z6PBKl3ObcHqWaZmXX2eTC3N2P
uR/bbmrpvzsZAKrqHVV8w5qWXCop8XsSX2p9jDeouZnl9+OfOlWhwaMQJhnny9VTizINjiTR2ula
dfhIrfetuexbiXvDTlAcTM3l2Lw2V2ofoXef3QPTGj5allcu118d6u5JiQcmXx4psatDf1iUnXhj
XryAyKDFA8zyvBJyQD9jdcVJEe3H0EHNaNgE7io6lnO28ucHG1f2p1RQz3dXKoWzFT2NRj9rquUB
Pw3nTVJwhi7FXUdQbiCckTbgEJAwPH+tprSbRhoZjJVOigqPlZy1kDyncikjzVBPQo0q5NAndPbW
ueIknbyHuAERWclp3ja72bJVHFSucYQmrovNe4f2yKdd1bntgtjk29TgyN7erb91kIPW8PER7BFh
8v86uSmjZfxH2IzWiXO35V0qdPTwFb3HaIxQ0C9N3Hc4FWK+FI6Lj3U33Eop3zm6u+O4XErdi12q
1KCGM10cMjPYJOZMG8knzMAZXxuxu1ZMRzen0rFgE3HCs83rU7zsOiLTHg4UUHILcZXGSQBMU5Of
c7w7siHAP+SJaYe7O17OGS9H4dcGxmBH/qsL91cH3eRhxyUWk3fSg9W4RObxmINSAXB3/mur7ppy
NAiVESg0Nx5rf74uExDf+iRWQUMDKEFjZEl4czGREtPB+B3puOTa5iUDa4NbbjhAnIxsqoTrY/y7
fcnq+e+ksJFS6DOXDzRpqev3Ck/qsrWXZK9HjyX8C3wd4t+sQYCDOveD8F8NQbxSLY7W7oowkb1p
gONiG00Qra3DRyhMxtqId0CsHl/cycQWO891rVWF2P03RmJhYlS1aBrTj5Sk+A/MNFz3lNzW7hIH
hqahp2Rs+lw1cCVr3ZqWiNaugCbcE2rlxgQmvkrEfHmzKFKzIVhZziB3HXueRc6x5wrMYUrztPvW
P1D1ricuUTGzPDpFXJjCwKDHlhpWvb1WctY+L4b+FyhExz7vESJKmcH6zj2uRp+CrY7NhWWwGZHC
bLy5Y26ezpwsDxtHpPJBVmjG2RnO2dAzUD76sbSBLPk19HkIq7guoyddSVSKXUNmv9AF3e5ke1op
FTGL8VT0f2c/lrCcqnsb3/stFAjzJEPIvTUZVhpC+CIjXQGwf1M+LKOpp9irpCh0tVKUZffkO4bc
I89arWuJIZvRiiHTdHAExZDgv59yEd+TZuSvZFz4k6Svo+IVbkB4oZtwwRnBj6AoztXJMwgLhXno
C/nzWvSHjtYLZDBM1GeAd9YuocA1xebVV6hQXqEAuusgMfi4IyevwG/lgDSkt6PXDHnE2JsJr/CM
7d8GN5OOJ8zXWf0SIItnBip9EngTog8B5CmjW3sA6ewuzuBGTWhaDFe07zaiquFOJdnSFcWcD6RJ
AIFoLWpAX5zsd7YRClZYlaguWcAYcZXVBpXuOa5p9bqZOjpQZSNiO30/p+qjZhK1G9oUCThKFPUv
Kx+A6PY+pXoYRrpwGbVXR58fVCGg+lIVif21OrrRIxQ4xxHgvlHxNjrNYMQhv8fSk6zjh0ZwhxGg
MOMBfFpvXLjry00N1AwFX8yCO/5azHRcbDn783NRhqbSrxz+5AlPxDhcIqZRgKHQx6TNyGsIw0Gf
2cMMynV52ddZRQN41S1KiNj/FhKgmAj5qXOpWc0uh1CZMe2U301FJ4LB0EjbSIJsgJVATISYfqJf
/G5e6E66oYeLiogxODEN2VHNy89dfBR6BlrQmFHjd2TRIkIZepcR2WJzwUlSze4V6ecqslZcBlM/
mlrBSGncTDOdufQwtd+kj4ajR+CZeYSc0xdegj+MnB+hM/7nvjdalmgKQ6cMhAMD7myFZFbkk26q
7AsRQ47T/dLZXbhgi4nkB3hVg7zzye3K1EOVKe0rn21ilq5lNdBojFm7whuFCKxQg4XSY2VAazH0
d6xE5lgZu30wvy3DHSgvXGthoZQqaEz9xv6EruneuyW5www4n7tLBANbZqEnP+uaYQh23OzrSnT1
rQDZzH5BBClHrQUlIAIy94bDJa3751M46aKZF7Oae99YrcJhe5SSyW7AL3dGTyX/NtiZE7Rjr2dv
n2wkzkAYWj7lJ6OXIU2RbF8Jxp56gcGJepQAs/fqvIU56c+1jIy9kfy7LOCXsGqahxcmD/vS4JdH
WpVZs2w5KFHAXffbiGPpcmJ3KtqxYNoCv1KQ+uHhuksATOna0RX3sRctdwNHlOufqBs8utjWSZJF
/4OSxgPu+W8pgSLIL0NQvA1NN1mBfode6ypEGd/21EeY8KiRGNWJSHQ/WvQl7glMswr0Zvg8XgHV
r71X+nY4i5DHuIzsf+fDkoViRZeBUdQLbpaLRfEvMMxbouoYLLXIwUQBCHmhsDLNHcNE2j38YdZG
4ipt/GtXx2LctwI32Um+gyY0va1fCloCYXS4nQBNqQ/UX1CB8z7DgO8cd34zPOx671qcoZH4glwt
bcuMZHKlvFhtkssSLjrJ8by+wAoKyrt1u2F0bbafK9KaaUPTvDz+eE/vpdbKAPqMD2slIUvRX+xT
X2tAWo1JBfaBzjcRlHFGZ1SJ277K5gl7m3ZGLGdk+SkbV4oIw5wGEh8CLe5h0SL0mhGffejKHuja
R+WM5gUr87Jfpf9BgIvlked0CoA8XKSLmatzuqWHUjukWsZ0LdKEXRaOw8SeR5w8ddFrEywhrcdd
isKwgPgCm1FjWKHlF9PF15k/YRvkwFc2XNhfk7Eb2aNUNiPULmuFpLa3GFWZHdrudTtavtM1t8Bv
ScOZjzJK8rbMu1qfZMK4P5awIMnyv/3j+lDlv6Waw/Jw9sL9BPhDhu6Tp7LWDqbsaad+kaBBP+nn
Gh6B0L7QoAc6XVm0plnJL8r2vX8uQXvb4ta9vdxGRpKpdwfps3tf7KxQGvf0kuDvZZ2f0JG8z1GQ
aBTQIjff/FE17JkE++Hq6C/5jOFPpGVP8Tc9mY7dlT53Tf2tlYMZ47r2cCLJnI3mvxeOAiQyjhWg
7WgUv9zjRf3OeVqXTl9YSRvoQED9VVds3OcjKy+hyK7HNdbHch1Px6G4tLcLSnCOftyJRHNvLTLA
/EdenoIPJ0wVZvJR6JvTQ8sdFJnBESRLRFk2+ArsYXYEwDGQEbpd4LiidMrKb3At9RpXwqo6hNPq
8/6//qibfnoZGCGxkoecn4jXBL88ztGvBHJz6395oSg0TL6sF0l7xPOPC+4CRB10UkqPwIJbGlQI
GhAk02bS0bUHzP09AfiEDfrTzkyQJQL54nnHGlhqvNkwy/QPAIn2q8YRBJwEOPwLCtHOX97YqHyK
DmlYbRJhGb+AaBf0C5KZgIsEiU2E/2ChhLtVamtMWllcAbxHZLs3T+uwZr2hbetiWkK96XGiSGRz
a6RuvX/LW5N3P/OjCfgcDu2Vv7PZFL5xehKNTKovdh4mIPH4yMclPZctHaR8l4zNhkszlcHVi2xm
6u/PUn9wxRMLpvJ8ul7h1wJpDgAF8lRuJjsmLyB0XggG4qzZ5ZsXzWlqWX/2Q22w6wxJ1jA1ueFa
Mr9jr0idpahmjSEljVnQA7X0YJYVzV5SZHiyLhueNoxQa66nZFsy73cmk4ndkdy5Vm2mgH0xq7VP
6nk0PP/Orx9MpDsKHsWoCe9pKqqM83sqM0wPV3tm6zACvdabPsWsYrzb5rCRbSWR0O+F3F+14ZVh
0kVKSDVqoz/9rHOrl5rcAtdeJAL/ckI5bn/JrcCBonw4pNcfO/4pWUoTB912SElJju5MDVpe6IKd
3CU9py0DjfAluFKaCCtCVk/L8yH2aq8jxa6iEZ8igMGmif+/fzP24/Kd1M+y/slzEYqZBC++a+d6
KbjFLn5zRQCbbfQ7Rkq+ijVVfaZaXw+25yypvqZ1GkKvRktRZ66k6E7BlllJxcHAJbTtHR4LNyvf
bxg8qhSGAVIeYwsoiKNHl6tXlVpb9H2BdSvEnC22wVyCss0VbKJ8qLAsRps925+XCaPkWzuiE3KG
0pFXlrx8VF85bPBr3G7dW5cnsV/7+6vCgJ22v8RVtHTPSP287wOd7br4WMImKs2w7uVPv81s2KzJ
Ix2QjugjflU8tXHKABAHZkIIH10ujP/qD35i2MDHfVi1ve8Khsxn1ASwDcJMzFipd7+84F/udygd
V+KsBPdIiCu67BRZQNqjOM1p4s/9jpFVmHH9cGIIAp2hCvdXIQSkYXnOShS+XeAfgJeVNMSfxYzq
bsiBKXNyKxQuQYpvtQ8nYp6iCWRh7CuHehyKcxg1p6k9YkPPgT74L0layEZQj6u3eHkQByrzRv2W
+lvvfdPDS2l1ptowixPWLlGa5VEMOzjXVTqRd9+HkwoBByQ+vKLk+bDlt7YzRgLGbbRteUw6xjn/
7jC0UDI0ugr+9kAIRj0IhXBVD+jKwhb1sgnoVaWyNhXyhA/FT4ejsLw2o5lP4wZJboUr2ECXme5O
w2EXwFi2S6Gx8gPyBiUC7T2kJ7Q0InSDwvJ+V2KPYr3tvMapspfJQuPHe1Vm3hDn3GLAcVlQCdFI
7Lr3GQK/MC/DNwW51viP5TnBfjP+iLFCveuuAyjBb41Gdm24Gv7HSSvNsqKYbj1dIDCMtwetvpWY
SLBXZHRG+2lx/I4iB1+rL0uG2K83QVqmoTX46eoqsN+9rjcEpbjyTFC05f3k7/Yd63gm4Jxemw4C
vWY+1LBVUYiyuxt3vZTZ/ELnzdB2rlA+wg7Nb75zEcrZCLysHcgzZ/WQ1b+3PrSouBQ2NEMetwa9
8Q46NvKQPqHncvWPCM67vjBuVEFZj1FKdqj86sDt91hZcvSQhIhXtUgVx705V2URk4RZ9jPiyM5l
3cBrtAMqv7n05qnSIxsU4ig90qk7hG9B7VS9VBHL+338yePAOM0yxN7+SxgM+qArM2LZpelOefSA
Hug7K9mKFGpAZS/ix1+UdVzhjM2JCF6SNQqIlt3U2SnBWQL8dbVZrSybz8yNPa47R3yEfVLNMSOI
aVB5Nlb4bLlDXUZDs1RQnL9CH+MHsVo7uNmOyc2Xhg83L/zu8x7wcCe5tdWg0GHIXHC7G1yYFnOk
2tww6zp5Ao6rT2k7IUtjv1eqoOFwCjUxX/3a6laRRsQpS3th4H5UdxTPQe86yp7KQ0esDXh3pjVk
3ZRb02U5vOLGWdyR00ipV065aVi0e2nZBEBVLIPzQHEY6oW51yXv3SpRXO+HFG50qAM3bUEq6e68
P7Vf21OPJyCQImeLLinK7IjNELzLaIlRg3xxzPjMIHBNje4XeJcUOUr4Vhf++7K0SIhkBYVIEJ2r
eRuNpZOX9mAjRaK4QBDGGsD7ULnyp3qMlMNMLhXCQHFTR5k4BUZ4nd6o09hLZrEOptPAjlaPDp2X
OtgPWC7ie8pBF5nzbsMKnBN4+K46jgT7acq/PrJwBIlU3MGxPp3dk8fstgrApk2okEGG0VydkOL7
b64HawCxJ3i/hWODeSLIFUF72KK1Vs19d7lfZjpIBRFaMyzGuyMUDAO5iH0IekD3RHSA3W26e/U0
Y6zpj721yMgV6L/ZpSRWMS+t30yOw+JgEHUR2I1h3yv5xrBNpX8UpYUQNKuObCnDLrEbw7QW8m03
43DIiLIMTRQ2BKLzQnASoj5NguNRI6T7mYM5aUTMZ+MSpjpXZsQ4yIN02t8HAdWUVaD0wKD/xHPI
++SoMuZd8gqRsArrdo0XocLisgf2IzfptEpNdcLxzhDCH2R2AOUcmFIuaFoXbNBn/8mdrEED6RSE
git6Z+EdGCUPe9EMAdiwkYNuA2PO+5fZ2Hc3fgXSsbsVlM2D7PX7IJK7tqk6G/EAuhs5WNKBa0Fp
tziqlM7EonI2zOdDLfGfK7AyBfaod1c6uMlXL5PfMN+XnqRRdYSO6nGKku+S/6Y/0fpGyaFuElEa
ZvjaRXejuhv0cCnChVAP5cuXL2zr0/y1ovmcB5pDzUdUfIenyy3t9EIr+pdjfvcc6ibBu9tg5iF/
3kJQ1x/Qj9iJXsxTyBFFNXo66FavjcnFcrDV6P9k+9ACrA3EImNVjgMLcpvUf9J1eHvE6UrrTwN3
F3SQKxZm4QeA3W4XTq7rat+6R22R1T4HtaT37BRaNVpvKgHR23ELzAuIXb1D+MisCMHD60nKsACQ
1+VaCiyXCSdeyAFWwy/RmHntkrPmDMcvek/POPkcaFelit3WgaY8rRItoKvqO7EGko6S/WzWbCll
d1spR0eNt5K1wThgM61fjlyOaNzCxEbgYkaDTWQwL3f1XuaaTwHrs+ltjAQTTUdUzzLArDKyfzPC
Ns4eL+2/oaKKSbEZjxP4yJgSfn8rtIPfn5y1mL3HRykDIl5OPmDi9NhcIa3Z1ow/yG4J1RF1U+Ju
QkQUi1TVD3L4KPFW7Kva3Kv0wx2UO1ZRtX+IiJDMwWThn7iJedVNNemLxa+LdLU7LlwpLoJkxd2p
psHiJp8/qQkuEeE6JnpoD13FngABKCTYqThu6EQFxNnJHLDjUggfavi5mobZgt9MRO6JGzN7QJZ7
l9G9ALn0lKSqV6msYXwqXKOPHDjExoNKgLeCyZLyheC8mbuCfJ3zE6T8EKWogFKUR0PfxZXXWGlr
QP2S5CR8DpJ90gZgn4xGqG+FQPHi4gxKrD56SyeqDftW6SqXtPqmTyJlEG2AqDJSEV9izZ6saR1S
BAtrKcCxYGr0PYB+VhQNXACjmqoMQl2kAuh20QDV0WdjDMigwtkNlykDw9YhsMq7cy7+W9e6pv/p
f3aSOJpM1Iyy27LeiiDM8HQmOQ7sv2gvNX2DRS1n+q9YAXqk1b0ax/75VOqaYJdh3nVEOUhGkr1L
OCT3BgXl1/TgQmrgNJMGS7j1rc/+WZPxs7iMcZCQgDXxRsta7larfUsyjkXafddjpeP5zu9r2u2E
3FBUEp64wtadiw2iXqd/DbIeOwJpz5vBHyiqTmc7//24Lf2H5v3YYzKu872HEiWMFR5II6j5XxkV
oDne7Z/BLgiZHrXHTpnySKu7JB5kzVHjqskzC4V4EuVfKy7f9JIeg9uJnXHkObvHaSKOo0EE11Pq
MhXmeiTOWeK5EX6wING6JJJPyy0Ku30FS1uey3sIevunObltc6hmt7O6OlalEqVsjoUDAnvyMkoG
8Us/Mcq7w+Bk4qFX3sSvlbyYBDKUyrE2RMIz62tMeI/HmbpeNLHQEMViC9L5DbnNJBJn3bHhzI0K
FIY63zMLJ8QvY0lCIpa2pbS1U/4vyZyIpCEzH9b/qBeDjm94HV/LUrHW8qxvoZW+xNnP1YHps9LC
n1+GacJiGfhw4PFpUzV+PYI23hOHNuge8tbRi1bq+poBU+PYY3Rst92421JFkgxpRQImUiQ4ifkg
Zdzy1eU7vHnfAPpxq42ubklT0FqpWxtoNFkcGPv9mfe7B9Ip5ky86Umd1Ai5l+UU2tVCTOmFOese
rJ+HImCGsYsDHdeqYTDxyo7zmTYBh/5pvcCi4b9hSCAVuH7g/CZ3P4UFipyr65Uz42/d8PHewprJ
XBN+duwlfroIi6mFDCboFlMUbs5mV050ts5sD2qaM+J4WtucdiTJkrTKyH/KgjgOIcx6/JC09e8J
jHYJM7pw2wKHmfaH9yOlmMHzdH8hNwHgHAie5nDBifv87ztP7taZT49FIdjMGiqnOf7hqB0nA9JS
uSgUmzTau1jtRxmp1a/dKYI05a+8FKIC6qFz1DNgg0TXgL2d8hFPp62m2+I51m9kJWpfPtUVcZmz
cv43UtJ5bccreYs1esfnSk+VzkATOvgdyjXXraRXEF9xyUZjDjC1BW/laO2c7yLJepTfLO70DZ7x
lS/73sQYq8+rq7d3qlBGRBNXR3oc94vFIAVUiW4WkTHf8PTGyQFKrlYnt3tFjhxCSQX2L9v+YRQp
6U0Bow9piCdICfEhmQibRKjdN8cydK9npykz8MaMTj4vC31Uf9gnjYJtRHLymf7vIx3EyzcbIt4m
MVyeaxKigCsf7opgiO3GPlB3yxZlLEo3Oa6hM4wvqglxlYsBAJDTn4GOVLXx8TzAfwlzwoztUYQw
rxmVs657oex/O5uuwikyhlDyeK5Kd1k7tdoWs7LYa/VEISCK8N4m/vVFnh/yMsHbVYGc7Bsk5LCz
Q/t0QkO9G7JOvJO7h6e8lrKJa/XWVEFPtx64MrqK8MAoRe1/1ZqSh/oN5h3rdmeApZ7glQbXxL3x
1qRA2YnJSd7U/YJIgv1KmzwBQf2qLnosWIzpvhFBGMQXUhxqzG5wjvqqaXebmEz847eYTS4mqY+N
6RPRZ2D/STLt2vTJDMMSIXLBPgpcY2mAPlqiJWM0o8zQCtfIPvrucanCcei0MaYjkhanNP/pG6A5
7AJ+tK3/Wz13HS5td8HlZC4mjA9y+kvTwKEvHD7jVPKe2KSH5VEp2sbNVA1pUqZGctxRJXCsYuWX
YBTANanaGSS6YV8BnFLB53xoz+8UeCaoazhbWIwYEjQ+7spTtRZgLrGvgYDzEICUjZ0DNTuJxueY
52ZDniNm95TwXIKqfT7hO7nncnANYVyWSH5tS3LzUt/cPJUlXBlyGAxM2gTR5hUY6isBHO4UrMzW
LhNGknpKqa8rl8NrAyo8wWT9JA1jXEDfDTu9qankoiV6BoEB0iY4z3EH2JvHcANGAxLCjNmWWFpI
nA54oiAn7S626zwwnfkOMwpUPiyLVIVBYbLOQhmxhEj8ZFhCZJu7dhEmNwe0dxF3seYcTG7oWExK
VuT+4tfOzKrEMGocmWfkQ9kspGi4uYjtfp1HEtkb23+QmmwfMbW4Jsp9/ZISNc82jlslzRLO7Lhi
r88EGVzbH2eXKAJ2aTuu5139XFqgNGOdI47SBvuWD8NLje9rMl8hey3z40tJivatiPwtzW42jg+w
pbU5L9fZBhQWjtjQJTFLSUpKC7yYS2mzCzts0RLb5w6FgKE/JYuflD5LGUkuXKl6qA80bNFaMy4S
cR/SUQyMngpRLX+f0r8WK2rmBZaphppfEBPdfnJaoAMbBKEQjRTkDmcwHCvyMSWFp8Jpv24qZI1e
4jq4CXWlrbklVcOWkXQZDugq2mfLnEluu+aUN0r8KV6mZ+6egB5mWTg0DXVMAy3XfxeFsJeg72L0
61bOd2M1oona3RY82nQRIzCzQDpWkpwLkbaKWWa58s4iIPXBLixOjKkPg/KZ5tvM1NnHfC8sZ9UH
b0vpCveaGza60KoZc5jorVsDVy2jQCdg4FH2zO+lwRZ8zdldojQIO0Giy/16RiUROpWmyEUmaI+j
Vf6QTGx8sLMPrXpK2708yyuw6QR1bnB7c39nURI0iDcj5QjPWnoBgT5ieByHnmRnEiz5+Y6CejrK
eroIlTkKMuNhrSpEwP+QnTVaAEkN+OKdKumLQLzvSdPTJSgAflUR6ZgDtfEcyFF3v8nBz209yAM5
IdXhZB1ACrJc/T20S78OJJRimjJVpkPzuroPJcGMVqeFBZ6dwu97wYn41juGkfo27MHAm127fKGh
62Dr45aGWqMvsZExfgnNhaNOu8ZTz7CWrNnyMG8+UbDg0dcbncJ9Os93EA9bm1DFXDWSvM5a21yc
QJxJZlQkX7aPawLsakL+1iJPlPuBl3oaTHoIbJbud5Ha7GP80fPmNmuFqa2J0CEltzhW0eYCCJFM
oyoOFdvVcdUpDJdztfMnxZS7oT9Dn62z2+JNTpng2JVO9ybChf9VLz34wAzYUJTe2Upfj41UG4tI
ejMXPHGGJrF232pe8ZuuzzeqPUIxQ6gM0+EsoktfkRdb2xa2raxY6refVHm8twgE1TUPPh5386o8
IFl6p0i24pO7ZHb5DdFEHULexPt1lm6ZFH+BPw77CtAJn72pKYniMBKq7uBFOGzcdmjIaHViaQ48
DfStdIyNKEyEHlsMbp32+gOG89t34oDN5LWAEpYEM6do/dH17Eaurph6plxgODar/G/xMK7VE/GZ
z9zhXdxWnXBZcHPzEUujWF4xJsEL1/y4I0LeSWbmSaMRXvGNZxws0xIgy3Xri5jfGe5hnkIazdz2
cTYFMSCiFW0fGDBAEwQhGJy9sz12HB+zmbgOvpgy7lyoPWxkx0PNC+08xWaf1uu2d93/ECh4eXzG
wUIEbD//T+fXInFeWLVsDIkYWgBEOYNoNlQzo27/Dj9PMWj/8WBKf8Z/64L5rgnsFUjnNcWQ17/i
BH6z1NiSoIy3XWDYUfIDsIPskBvAieRJT85s+ALxJzhNRpZ1Ogpcprr5RmbIuInXILMjubsSyB8Y
+x6/haK4FrdDJwB8KtTrCVKgnF71IfraASsXVEzXe8RhADRPICj+FVfbPlIWgWncGVZKj4aQsuxG
Q8k3e/6l97LNsWQT9RclFnNqvG0LLv94pofPtaj4X7ZNo1xo1x3b8sqLfCm4gxSYVMtrseRXLnuB
H5g9WwTDdEkh1aVZzdfakb3sMI2NLCX+zB0wefJmRv48bLT0s5bleGCVEMR8J2aeOl5z52D6QWFk
Kv/sVLkObQeDeOwXhI3e6NGhkzo25RRYKJbTWHe7M4FV60c7Zzh1fE02+H/4VYPaSdLWLZ5mtgf1
ZLZ2ngY45gnEbz5qkQ/Hbv1Pptg5IRbYmwMz2y+UmJjedGCSxmRYj457eS2eP4VJe+BKAZiOzNoc
+YJGMaZslYCdBgfC3A4fVN7Hk2jUz9gk5wsSVTsBX6LQ+EjtO/D5DPuOoT7p4BezAgfbKwItXBs5
V/KukWtX/mOzC6rdpLBXOkmeZqYDspUo8Ng1Oie4xO0t0YDBLoCgPSeP2ivUoZ8GxyCvPJpB4dBc
Lr7Lf+NQekr1JL0Zek4t7XuLtC06m7T6kd2uZynuaMrDNKHuX1e7p/UgTWLm7EQJK/NUJH2hzEqE
2EeIg2fTAIT1VVf/E5Nu1WBZdznIKuqGhx/DQ9VrPEqjd8OZRyVAeTcKvs8Npw/FRVFk9j9q4qrY
aafxQgcdd+mYSsPsliP02djhK0sN+6Nui5or6hzONDfTGWyGWIb0sM43aGbydFIMEmURnWgElTUI
r7kU3S+si6eql4Zbcf39GmxcB8cL7P7+y0tzMNgb8i9ql6d3Q3D+EHvtNud63E4aIMY26Ru3Mv8H
xU8WaQik75bX8xjSbEIamIOi8PRYW3J2XHhsWwk4sZDP/kHWvQqnHgby5ybCMlcE0skOBlpgZJV0
by7VViOR5D/sUOx0sFi9QOp4OYT80B5Ly/UK5r3r6VJfLJoaGBFJ+wYkuy+K5b/K/2ONg3NlaPhI
4rodsSQ7uBY39dMewDUXjB83DtSquut7OKgZEsE/EQTaXheIBe8cLIKTcrjoSwnOoljkaGKkcAAS
yZx1iTOkJYoDZNcOyfqPjkzYi+0O0BvZhE5ikxwr1wk1EyYvJbEs3COGZfulxJ/JN6OURSBpQWnE
vveVtLaWUxGMs7QUzm4ZjZeESOThYShLsNzi6HJCUsTkHL5yN6Di7sbwfapBHCmddpVCF6hEuBeo
lwjXeJ+SUx/vPKp/AOiC6S3lkRt1b3rRHfSsdHvQT6+Dgq+RlIq+g7vfZx6vzo8ssegIZQIU8LSJ
XhkBVX883kzfBXBkrsjE1UrBtW4EW9Gt1CIRaWIbbBPGbws2RzMk2Vw8I2oBPa51eHVkEjazAkOU
ZwSILSKMK+/rgeAwmBTIPXTs68jm1cq3BbMOZl508xxCFk7s0tsDqt6Uoxcqrwg2APRE0EZ8vN9u
I0JHoMf7LIjyANuMRHMXMn7A++E7tgj1e4aMnGmPcnzT3fZyJ6UVzZOdaMDPRqHDbmE63EATVZyG
65RREuLHScJZMUg7t1rtWw9qpyjL9hIA3OU3xy8n6XK0LQsvHKRMGq2piFFYyPnNP+g0P+jEUDyR
Zu41UYkIQuKNgqCxj//SX0a8VnsdCmeIkB6rw0IErO/j//MGIdWFU/oPHTtZiK/y1mkLb33H8yn3
uhpV+sQeFTZorx+gG6n7NI4YvaGgVipHJYajupcsKe0dWEdwm5yNbJmjCoVUJxeJyWxdGS0vpLPV
kCFZm9Sbry3CfaN3AVvPWu5DGT0/+OFu/XOf6F0wdq2CezPj/t79NDH8Am3TSBh6lxiklZ8dpV2X
Fkuze1O9veVI9mucgEc/Xn38AlPF4JZenaFVC+tRRjRw8b+Cr7InHsI5Vtbh9v9kRTPQMj39i3Zz
ORaR0IsdJKDso22kfrcveL5RrDdGeFzwsEaG2B7h5g5/JQKYDo5+2PVyXEYEBkC11rlc6V25q3Vp
YT/k62PCVyO25WJYcdrQRFaVGY93VpSJ0opwcmK2FuQa/5+77ten7cMHA9F1kSGorw7m2YCozM5w
OjlBPjN1H/bLwVgP6AgvE1AfWobKpXWevIGsl4oVjTcZIEfqpep+8R0VeWUg9PYPBN5JJgrx77TP
4/NcUvAbCooUXVTwNpPutKRjlgavd2ldyPPBh6kAX8QpYXneJbW6UBL9YNVCfaIsmwb6O59pABCU
Q5ty7WK02EqtD5YfOYbkCtTMzwQyX99kNFtvr12Gx4c9R0YDXQOTq9/v4CN1i+XJ/GhdQOOZ6aTs
Y3lG9z8ZzteuiaTrJWafYuezoO9emNOOE82nM22lpMiU/+MAEZtDR3tKzFis4Q5ypf0QwuOVrs1W
YW4vEzPuiZc+cIyNv/ts0u4wMAG+GpAFc8+Y1yTVuzMUXu0MRBaGMEFSQhcuPLze95bxWx/Tfxaq
E/EO5S5ph2pkA9YkrV5AMQOI6YEDKOA93nwtar0Jt5MXI/LKhYej8kFtHGXZ0XMOd3FJmj2fYMVo
v0Mu0C+BgmGDhEM6AUF0I7Q0fx6ov7PVsV98JnHDmBU60ZI9PUFWv+sKjRHhKtn75YR5MQWQIW9X
glT4OoSkJ4CoOq7JLGMNBnPqr99ZAXH34zgJ3/waJ6AhblXryNcBFGJ+mbKuCQA7SQYUip/vdI0n
IRcI/xMEWWREW4JHO/hL+e6hZlo3S5XPhcMrBsFx8A1p2dC4lMB0IavETmZnwbY1neP+YwbpJWFb
DLpubl05A06djJ+yQ9zlLeDz97VrZAWsq3/BOXceieLwBq0+mhmepOUEkY/LbXR231atBqcQQwc3
bR3qzPazgYg7juTEePHSTjQisr+qPQdD9sUJqctfHc03EyihEcHMAl6MG5qB0McaEJ2lCEU62TWZ
oBlnb7u+AKpSWJxItq1+jtw9i3ng3jSRUOkdtPgzGDWLX+EdX29yzgQJkpSNigX422ji+mJkeHXK
tTFEl5s7WmaCyxOYw5tUEdoDNUKqwCDI8x1v/KeZMg5+YDDif/ZojNV+qTIkYHVKevPLESYPABHW
sSoWoCnhQFVH8trkHj946Q/gIRq7JEwgnbNDKod/J6BDlUO9va6FMlOhWgpvHgDDjlYmXGtqEkeC
bsudjQXg1/K0f3XP8RkqjBpIQbwaJmtcfa3p5KzjRvH94d3dM6EfCWNQIvgP9IXrjMd5otFZL7pF
S/nn8nBfjEffl7V+NUBOR8F9y8BSI3eTmR9jWTyHZ+y9HfUMZYRNKJrllN05AyT3fNxsgkTkhBTK
V5fLtUvvKbErRrsCYySs92N8jxBiHkZLUdhltw9xCzrU9cCAz9mUXtVGhJrVzZNiml1t+ohxz61V
k0pXYv7LdyOTxMKvfhyYqU1i0ZnFsYThsM/B2fiGvBoHOm7BZWwZfaKlU+nBTmzB4mcIUPJQEchg
AVSez8ML461mLxF+jHrcCq9cH7Wb5vAgMMjLMqjOlhwzdaf4cEfB/XUCqSzKvLBUNVajhXavIY4r
aQWtD7PpBeaUhNWcpZOb8AC4t1Itz7Mw/OCw44vHN0c4Cd7Iiq7Pd1ZYlSbDF9oNJZsi2R4ObHbN
4uZe5ZBmUuklo96acsp5gOD5heJB7bMJU7lvByRsHstGCS7+bYvm75fBZEpEbIUvOEx4YOEJEnOx
Q+AZrEzhBAJT3ZxTbnYI/Wl1vdbrn3EQ7Rkt6bQ5aOXPDp88L9qwUrXXDzPXQOsbKbpjXfJZZAz3
EgpguNBRyPdyRDgs+/KuqGA8DG4NZijg/KeshtSO1Zmj1oUGqdp57r5ZNwoDGxGj4UQoWDInCUbG
oqs5NDx1v9Upl+xNxfY7BwpIR+4Ey4+A2Xx8KP7rE64HPfxBAI7AFtkjobRQoyb7DVazdsrahS7O
hdNGVz1HkwvMFnvdhYsrFde6p2SLktUhS0lXWPSOIVZQTuiJ+EHbuCetwpANk9SE4Vc1jXOE9vrh
VVnbG7pJlSNXhcqIuV7dcI5A76VNKQ/jox2mHBeAA4dDFW9XJf1xbE8iBgt9mBzN53M+EIdfI1op
irkh1xOAN/7zl63Ap9mUfN37FFrJeP4hIuEilHpQKaR6oBzeBSJOMMuZ6IUTOVG1qXmJjQCX1FB0
CIz5gPc94XhqM0zj7wpk3BtLy+gXlAjzpialnbaDveqt0sBWGiLHsOjfyHp9VPTuTsq3vmn4D5/7
0HQOGli5l4nBWlv4HdoE4B5EbbBW35HO5/bcHjU9mqR7VqEkfGHAvOUkVcrvROv956oGHcogoHTU
O8JkwLuqeF+lrh1losL5TVCd+Yduli3YW+3kenHe8XvgG2JoXzLhsm/HzzrkPWpEYnagPXyfIQj8
mSkfeqFuQqhkF3G2q/E+7E9w+/ETXqo/QMB+ufDfHPlQSEcf7nS2DMVfJB2S7/kcdB+e8BubYI6G
j+LWwKzJ104uQqC852fjPV48+ExZZiblYqYqyhf+y8OA7ytRtFPsDWPGHh9S8284ZFE+CkgJ6hew
1Zf9J0oQFBCTd4N2civoDhuk1ucR3CwDkeVbQgZE0cPsvHhMejSJ7tLnTe+6FVjp3kx5+1r/N4O8
jlqtfhEC46C4Vx2ry0JV9d9vn2wwoKSgAf2VMr+9fzESb8kko4z4qUqrFdvIgPA5mhWTfuQHE49+
SD+4RLmp51JQeJIDOQJhCy5qzz8stT+VsP/ygAnfhVCB9TdjlESn2TMnTux6hLgb65OkRjYlLjIp
FltyR+DlpnarvdE/Yfk1Gay5Q0v1cLSEoJkb2H605fcmRLvl7vJ6g6Tqw+WPEXtqFh6iUNOMiynb
Qhq37r/XK5OKRdBERL3modqNtH0PA8AMk3eaR+XJPeu/JyYl083khsJorYzC4iVd+TDlELzKCsy1
zQZQRrGi/JcNzSAeUkaDtnoAoHXjv3Jxx+O64MhDzppxHQh/NfYzu2QnuRMagSduO1LZxhLQs7J2
fK5WaRlC+NnYq/lh0Q38bg2MKbS1vpBZL0iqpEZdJguddiE/TBC4ctAHGYj/empSDwHqAYjIQfEQ
i0eYWqzZ40rHmsHv18YahHitHbDWmsiAOlpfnOJUxcf0hweaeCAY9LFIGeFjfzVZHLrxiStp25Ar
evEesqxUOB2D8CBeU2Pu9UIrNP6iHhwGzsJrmSBbmAoxfdAdqZJTnEzbQm3N1HrPE/iflB72AaO8
qDaNJ4cxVwED6Kyn8vYsiF28We8eEov1B00GJKUdmSOP1mMPJyc2MZFMMY1547iu6qvGiQZcQKAl
EpzhmNljm3M+gwd5Pio/tnJJdPftvzIwxTjr48moTRj0uhEB1FV74pEIvhHzxGyiQDu4lihWqsVY
rl6p2vZb1aPelna4mmnrGc/2Gi1zMVuPIX8VHHjKa0Lp5Pr1x7cfMAv1ypcnyyiOQ9wVpafW+7ap
GHmKsfG7omj8GiQYhzVnKgMzN5Q0UjK8ytseBcmk9ukUSP4uDYqlW82vkxYvB+GYgpEhrmAbN8Ag
9AnsdGWlR0sikX7FkEl+JvxlBvjq56mrGU/0T1FTcBvLPG81lzZrYkqvzMFahTlfQnNosXpIwZK+
WeLl63thMNJdueGFlA9y7lY8zpepz05kNQu4si1u1nfBWC9uhu5a9nDEP2sov+2DpWlnwB47M/KT
p76mJJmdWT6pnHI19i51GZ9EV5BeezpNqu/oUANv7soXceUlh/b0PgrhokwHecCffE3xEQ/hhlv4
jPpP0dC6ikB3HZrBhUDq3rwPzXFQwHEpYcAxINamiNyJtUH5B+3wMDpXs1vQ9N3kLLI9NLPp3mS/
XiGYF+nWIpv1dweCNhWTzSWSeHc41ATu784/LbKplKKQfMHiRbYARJb1UgJDSt3s57BGz/fbKzO2
VhO5bogvQOZ1eYR9fHcUgw1pR6HP3CQHTH8S5JOZEo9T1rVF7GVIM2klYMkorHTWkPJ/g/1NqbLw
m2s1N8On5ADJjlP+pr4zXjeHEe8jY4Rd3A8eOdPVVb6mQBwsWOZkZ7Y5oFB+1JzBaKKm94G/mx4J
B7q+N4vXhHBUks9pF85gdvLGIQjP1Q5arl0ZBe4eVEJYXenbW70/ohlZnAtKzgLQjVj44yVIec9u
gDYWHSJVu706wHhDogvhR6mJGDUdQumanptrBPCDkbBWcFQxgYG6V4DfABKrBE+01EDilJuOxBBJ
CBWrnoEkma5/EJ9U03hToZa28WtSY3bIMihPW4DDrmADPd/GepQ5zxGW5x7CPfgXQMWKLodJzhm6
DBRsXmZpjri5ub9Pq4FNdtETvYBsCD2grJA5rhuRIQgarEgrxhCOKBJz2pqOSz7Cskga/H3fln7a
vg4GGsO2l79Bta1Z19IjjCSG6yKy1xyE8QpO4JBD4+QMKh/PkO1BjVlipK+a+jdOzTEJDgtdSMSg
Ze3fxIlZcxkyGGmzNUgQa30gwAiZ8/TEqOlhTUsN55QlECtoxc9+acaLFKjWbuVbHnmfvRMU8m38
HoaMoxEiO562nOm0KkXouzfadmSwzxysA7WaRvbI6Jv3lIorp9hPgEKN527plV+lp6r+f6ZY7uT/
OCWtaFRVeKQvApMlB3f+tLGVELvz5H7cUsF0NpbCXtg3Z0ov4JmgN9QRM8/76seToI36NgfYYbxg
QtqnM2FM5bUfvdmm+VsoSjVTl0SS9czeYa1G0W1W0MFAUUs1WXQmRs51VD5TUYIlzd1WsNrX2KZw
jqlDOWckcYX+C4UBoQnW7h+N2cdVA4Sr35ka04PsFF0IUE56zNO/Lddw59Jm6Nk23EvrhUno3GvS
uOL6QELqB3XovclKPp4zU7zm+z7ufNxmj7waY0JnfiSOD2CM+/Pc2lCqtyOw3SQiVBEKZLR0hPR0
pcK5hWITDdnQaOVyXk8jQttUgK0LfM3KQTpY8TUxt77gQv7fze5HfRkrCUWYMsJCXY47mTKo3MxE
4Yj9uiNX3kkAQ2Gv8rGgRlBg7WZoqWpjrwkWdigJpdKXN7XQ4Mntd2DT5NoPBL5eoYdd2QkYSuQ0
V8GQiRPHnFXLXO8IDCXwpvWhomiIoKw4BppbDB/uoQcCHyjvsiOa2w3olMzceYTNdYYoKRmLTkBy
pRixuZIKXFeU/NbNBa9Tn28FcK4EppXVdT5ZA+KrkS7/iEZHCksV1PztYOa49rM/CwF8/0x8Tk/m
4eXcC5iUvm6KQZb7NqR3mMCTiBbWZwdDGJ3daj8HHtKAfoiBN6snamU1wS2NLf+uAOz3w0UdJk4y
plvxNg2lNMlozI3UazXDdcGssRPewCpHQSpUCz6B8DFp2wMdNrbnNi9TxE+s2AMTuC13e7KXz0i2
21p30d2zMjlz3yqLRJ8dAufSCJ5mAkW6wDHYXm++gvOqcSQLDFVpSre1ZYdLPbxph/B++3cJObyX
G93U+xecO/IYseKBliLyX+3Fl0xTOMPoSpnS/sLopXE+JW3a0ZocDUeUotD/cTFaHQNLH6mh7yyx
DeJ37un3XTck82O2LGKkF5z57sxhhJ/01KTJT6pMe6JkWfsc66MJ/VSCKOmQXK7XxePj0no5ZN3K
aOkJnm3Ghlppf1Cr8mBJoFWJcVXEjeNMKBPw2+X3x8phYbS4p8pMObKLyk5yS03yy8gpc/+xehtW
OJYuLlKB7gv9XOtTeQk3vVWsqyOtjjjlAA7Botp64vCilljzI2lfvjAan4gFi0s7C3nhkFjxWxLu
62TofNhVjYhzbalkF0lCXowVTu/APBQM4RmULVxI5pgTOo6Ti14rs5IrS2PpJ1A5QrQIPkzdr2zB
UN/2NB9uOynmFM9jekfjCkmvoJJLxlDjJ9h8YUc5M+1FWH53eOnb4wzZlR90AIgg2AoRDEoUFCcf
opF5RGjkB8WHcoufrMMGEHYCe1nbjZfsIpLpzaWpBasnX7k0wrmRWivpDWjvG0tt3wbxkNlqc2vl
WYGE3tzWm4+zROnh4HCwhFw3GSkvrg7yE96Ri66mUz7PTBhilyhU3vYTHhmQpVVrNqnBqAvPFsr4
0ifRGF9VfFHLkNHF+FlZ70MDDMC9loCg0VtIuwCIJK1SXzvjwoDGTtaSSop90d/gsL02jlmkddX4
aFlEc+gEHqdb2qSwDJGn4S6hKIQnJg4DMRnC+vip6ux+UNWXM/R2REzWoIKvgAGriNNENpwoFPdI
f2BeMyY+70KhMuAQPAYvCNkStRWGfGdkdkqF/w7HbZEzYDu6J+vd9GZjhapeS5TaSS2ENyLQMry4
hzXK749zPwpm9gAVbPDKh6ek5UjVNAl/J83vlJJyZRw1wuOUAyG7rOxUOJ4LKLh7aMq9dPmeLoJ1
4Zvlxj+4YbkwIODb8apHSToDi7B6wVt/ihXqGeU+QW1ZjjNzXdnj8SP2Z9ZrvdLpUlaLfsyemxEW
5q1OTnkkmVpuLIRjjzM9pkzRxXzKgZiacQCinxCs2wHuOpEW3UWSkFR98gHewJcWiUsa2FnGx245
NtamDH9O4N8xqQskBQsSrweBW2alBGoOH3moYaQkNzhOAB+GK0icZcJJQ7nWJ9qD8HdGw4YKyb08
4fYBMVdJFmLimXET2pHSI2t8Gl5S1e0pgahPSfkU7IYK+uGrDSIKnu2w3HK3RB5MwXmbCXH+48ca
8WgeTli9U4zE2zfz8XGrMpEKOpYUG743q91VBEB2A0rquAd5gBg4TkXd/o2dKbOt+DOwZYGLyEK9
l8VhYkNsl61N9NTaIg0ftcgC0NJaT3YU2duSWoz9jEhWecXFkLfYqkbbYzHNyIKZYiBoM/ny6vVc
O6fwYUqZXwvbLBJunKxCoIh6yAhOFpDvsU5KWnTzqEVml9qtoTa9zUm7sO6tiOFYU1fz3D9hLG8b
wHPNv4qVn0Hs0yJafy7YzSfFWyWZYlL2I7PRZcn7i2Tysj9QwyVaI7LMwxCxbK7Fo1zJcpxgtLMr
iuSGzxue2C/y/4/LdPXW1bfndWgZ52H9rqrvI285hEG5ke5peMeXGb2Giu64B3s1MM1H512d3i+X
8BxfkknDp6EblczoWXBStgwEUZZ+L6iseIjOe+/3LAGRiNzuf0vmo2jN1rYuSmDRCnhDTdH+O4+X
0NhDJDanNxrlXx1m6B4C7SH2PjvxqI9oLW9xWdfrCAjxIRO+Hlc2kqN+Hxf8tnJzwXpILUf4gYKe
+xby44RAtfqV4zgUeVOpwJPrNCzyE73sF5UyYOkA0Z3HIQyTWzQot4NUoZtNeEp803BEfWr0kdw6
szjnNipSvPpooTOkRB2E0yNK7L83LxOwvwikm7K48eJyBsno8wnr8d9EkV4RV4jzQzHfnXF7s8fA
d1Nm/qwTZxU8XqIu9ZzVeLcSCAn5st/fmB3vVfdPvNIxIyIq5PatkFrfy4AV7Gf8QL8CesaFM2iO
zIfsg2nSAlrok2QKHCv3SD6sAmAePuSeOp+eagZOqjBNs7cqQipspjDIIt9zttF5ZjtAdtWjPXLV
TAev+HSNejwQoIKj7Czd4mbibWCWo13YKFN3DDTpSZmPXsj+e6sONe7mlaG8RuoxW1a4qt9GJ3n8
93zo+5N6XnR0GXEdYzNndMZnyE/gxRXmViH1E606flRiBwzm7ck+/A5SfjWNFhSxUg1vvWdKt5jc
0zHcmAwPtNlo/cQmhr3Nv8mlCSITk+fRuAsaM0F/cWYHXsxDQDVzAFc53yC4ndAnOBikjEcwdAmJ
jLQD9/e9fkI1WNgt2fE8lyUHe3PfkDcLJXf4xeKkWl7J5qDhLhsVRJ2q1YmhNfctdd/IyeafsVIV
5SKVUd9fMR4mmzU/tccFPPOYdtnvRz5DXTI7BnCiHT+A4pKFbjPtlv/ldkyuOT43ww0Gb7K6hfcr
pUBMbHg5+6MyjvyRUxMOOjYtgaXsTSnS29idQoGtj1053DPbUltOWuBgg7S0X1/k5XJCspq54xOX
j/XZokvI6a2qjAdOaMwvK4Tnf/wfBFA4tIlIXnZnnRsn/udZYV8XlHS2Jz2omvKymXDWJHrjkJMN
IDRMzLrdEWWKTPgX12HTmIURKHt2FfSwzZvY8pP+ibkXEuHguWTelVYLTXLnZn8rVhymeyVBsLPQ
ut2HGhgqUoCJxx8Fo4BiyggRN7HeFmgIF8UW2tWovA3O3XRIZIzD38NW2o1IY0oassRgU7/rtgs0
WRcy2HyJQ8cYR2O8vnvuvo8dr/VEdR7cCWvF57z4a1Rc8/9dopnULRJURBt3iwSuv5UbPGowDGgg
zv+eYkaAVIyyH1OrnjTiKA0q2j4ukjb7t71MsJQGhOn1ATkzsUR/y+oeY9pZZ1KeeOBCA1I11HGe
fCfwOGVt352cEegiLbl9apHNT6/i52zAP0ozW3WIOG1Dhwlf3Ljp7Xpz2pGOAp7DoCJcl/lcL8w3
l54aLwY4vEbh97qb+rMTziX+lAp8pH4hAsljZyYFPllFMIogNUVnWf28b38n5P3loGbriF0vIxNN
NKH6cprqbJ8PtopsCrqk0cNP/G0fHCfr/4tNtw7J0nvcbpDNCmQwA1xHsD7ZEPQTlHD7CLxcG26o
pEHc8ep8vDalpobS4E9t9ltbYqWt347OlJNfYqy3lNrCPqFOgNAdD5xyRD9JyeKd5DoQik3E31v1
4D5rCTGUHEWXNfyTT5L1fnxtJhYFvJA4YDln6iG/pX3bFRd64a0WP48LNIddfjW2VKYD411Qem2k
ry3pfTd+tJ7powzdJUDIeupZ+ujtGsadq5MboBpHYVkkgEqtIZy/MhbQx8J52oRPMF0pUTbIf6mm
ImxjPTa6q1sGekdp1Fpw/rU/1msoW5KQpGQUjOMVCvn9Wrxg0rArtgdmNodtjVy2Wt0mRUAv1iTJ
xOPclHkJsrsRiOtCIJT9KGEGvQ45aar9t8lu/bKRP88shTytmbIJGGD8SuUPYCNEklD6SpcD7ZrC
yqbSI7Z9BJ0/IykejVV0LB+2J+XUgf5FqYUd/Qz1Uwq7r/jV3YHMknE1+w99q9JKPxt8YuNKXFfv
hiZfGBcmftoewIzS22zEaXIMw5Do+pptxNVqDtI5RMgXJj3je/tn47ivG4JNrkT9GBFE7YRbhuqq
HvDJhhlZmSoOJamhqgtUy0Uka2eqgOqjpsY+K1hJwJMPmTJ4hBxJWZ6fpG9yZAnzUrh6AnXewjiU
hJ9yQwCiBorBbuMQvaqo1d4FXXLFo+axCOeHHhyiP2CfPS9kMaH5UuF9noNIuL9ZeYEIaYlvtRb4
WdUnHrDSF+tDlGfCTnRZ6IUQ9GLHoXK2bknmYYsRIPrnWfa7AM8ZFQTeZGvgOJt15JObtRCSwAVU
o+5Yu+LVrHAXhbeJ25A8yHrWwEkJ5WzRxcIV/U+ZQG7emiXFuAAt46E9o6tzh+2WsysL+OZ1A04i
K4T53GqoP1WtFv8b9E2zfWUcAbmENcDIVSjYliq9cmGWBnIljEZX7UDDdvxgpUWOUWyNY9CLPB00
yIDFA2n0LXm98VxA5MLXOpGkg8zTENULLQTr3ROv6Js2MtWvQPuiLXPYvcI/a2XDad72S7g0uiHF
9WsG88lsKzexdO3ylhzjSp5Iw3PIIPVY76WnXh/pnvUgK2Xn3DdsFMOEo524cqu48SR/KKrnKTiw
/0ihAuITMuDU99mNKq6231Dl1fJDIg5tIHYB56mEtupHPPkGPDKvtvGz4A/ChxbOeNmFn4Q9ilks
iLBwStsBx80qctTvTS8qj6OUCLQ1D6NzaJbXNCYb9HbBsDHAe1NZ/dLXY/D4xj/+YrWFF1Pqjx8j
ELYcC+Vomske4ChGB4z9zIwDFoZbvMRX2HArgmiXUdfTK+YdUfu6K+4rb+yff7i4zKp3mqX0zYIE
yQcdwv0jNB1lrdH21G9dFQtC1yNFi62XiTvEz+v9A9i39Dh0jN1zmED11GIBi5u6tvr2vCGyb2gJ
TVITk9BrB3AikDt1Et5BRKgSUTGGzOXL3NwbLMn6leEmM+nOCSZgN2JRYwXRJ2QaDDSFGirmq2zX
4FGUcTl5xbh+L6vsxJC/9umB7wJ9BjQEMDjCw7sW8mse8Ybngm8/az4B0wBZk/lz10rBswGxif/I
RVjLNAeCQG+0MY/nFIPQ0H5VdS10QPW48dMnfsbiaQs/zLw0if2l+gbCBRJGgNLiVhyIRVAGSpNO
FI1uLVXDpuxGcw6H9g1qY/rsueBFpIXsMAAIH4G+Dtyi53rhCz950IfOinTioljjwK5J4lDETtGl
+v5BYtwrNo4Gnh4YA2k/Ka3v4HZc+F7ju736U1ekDg40rV5viENdWcyMgMlDaDo4EWf6biHRtUpa
nxe5Oqszb3EguhFU3aCd+qRgIoVc9oGmevHuTbg9zj1mr9HKOVvB1ZlBhXF1z4xlN1kBj12Yn2HD
ASNcazuS9P8jgPu2I78N5d0iZVd7rFHqqIstERdu3H0dPAmxD6GcYEyK/tLoA39/rGebtJKFV6YH
Ef7hiv8JWlVCoF9KwdBeVHaGa497rmfipAteWMtnSc4bE8tJlw/Lin4xpB2PsZU4S/KHDE8WSz0+
LXs56WqFmHurXQLOxuMRoPECSrfiIbBrl/ZPcRIbMB8Ygb8MNvzqkos0wiPTQe8ZP9LHkKKdwC8s
lW0wrExsKwsc7qe0KkB8tKQcA5nOmEWdwBYRkY/bxaqcEM1YPvL0vUDWuO6fi107tKnOfIbaQg3l
VUNzNyPRTXVYM3nUeePUcFm0Xgjw89PbDEYIWbzkQmu2rl8HwCnN68RgjbcBPTq4pLL7FhXoXf2F
ZE2iQZ3YnOCXrnaTDG03l0MLoDDk6SQAljHnWCxyBMUU34qJaGFZQBiGKBsHf/HZ4wx4lcbk/Ykp
6SHg4cpg0ZMyNy79QPwifu6ITQwHvLqYZ/xgqlwyov3+tFhlfQzrYLJzb8rJMWzULJY7QMgR4DJG
nVn4x/fi1f2qQaqIFBw1EDvl0mzdVR3nX8qNb4J/TZm77iPF2v6SIqF0u4vh5pfsJsvlCi9tl6Vo
POwtdE1OCM1u/guZA+vOg3b5h8x7EyKvdaR7qmUTMWLf8LGSahWZikEfecbkZVZsElkDHeors+aD
5B60u8fjCW17GGaN+tSZcVboA8qqTRE0SrB4b4A4u04ESnxTFn9FTGRqHjuIVmBuNWeBAfsF9gys
eqEJE/HMgtzNm9Xv3U3Lh7owtzGN4+EpuS8XVVvierxWcPCjnO2c6cVuGmuApnxpmlEd+WkGzeso
ftYwrGEC4tjHeGBr9VM2gGXxxKfPWp3V6BIdN6TcU4KP9Kl/090tMJn9nUBq/Qj4u01bo8KvN3fR
+6ldP14k5AIiAvKcsQh0XhEffsPHp3ShApOb+SYzRidqnAb15zH9bsBTeC/ZMJcfAJvCcEThqdBM
SDZZa3t+940CvuxIcw4RGZnXdKsTy2wcIYIdImha6HICTI+w0JmAaAkZhzlj/CzgmomFS0uu2WZ4
xlSTGHlCJQUDvvV05ZSFwy3DUodECixJ0fQXWSEPw3yuaUhzpDJXsTQGwYUACYJ3DofK0x5L02PH
bJC3quuMMD+qRpQ7ryLfsFe/07qHZpx2nq+8UwP1i0LfZIHtDTv5Y3sEJSyZpRbuKoONbsc5NC7p
e7/i9gOUBovfmUUq82McMstw2OZOF/4Cwem81xP+FnGBqnpfYnx7u5ioq9n1Mng+teCKi2fdgV47
bOyypi7lSrQrMRD3YRV49aTjtqDCA5RKF9m2jO+5PmVWjie+cOkBTkO+Z9YFKSHLjxHDDafxQxsg
JpZeyV6wdwJwwPQADxHvWMtm3dId4A8oh2zd5leSXJ9NQ8GoER66IBzH5KcmWnWZCeOobJ0OUlwS
dHvyHaK8AQ/9LEVZ1V+izBkHuTUFOjxPVclo3h/0DxN0BBk80iGYI2Yii57FX+HNqnr2calKfg35
pv0/LACOHpbNkrTA9RefNcZn4bY4m2JLwASRKaUA3zRluJa8AtcLdO/rUGS5ucvObkHbHueDMUZo
7UoLQI2PLH+TI2IewisEz+4dRmgR1smQtWfUIe2vjVlkdo2VHVVc2hjvOgsRK+jtuHmOzv+z+uUT
fd4aLp9xt6rVfFPz0E0rl7vHV4KFC5eYfnGSi08I/rIF1ZmPByMzTTCfI0x/TTTsBMeV+K8FINBu
Of10KF8vlNMkWAdZSJMcy+gZEvnSfOOlFMMM88WQtNLAt4z/27QIM8ruQJ5nHo7o6wI3mczqdNMW
BVGzGeWCC5NvZ4UM0GwFBP9WkdhjPVu2mzMX4FleA2GRjAxuAWEVvI8XXPzNxtZykHLhVkPuqxkE
bPWpBjD+cQZinl17nf7Bvw+BEs573SDNpOkDKENwm4+wWZRk6vftufkQnFU+65o/A+ofn2B52zIm
1zPqnUW1IyU9nri44RnvMGhlbFNatiHFP/2o1AGiYYcazLfRPUoqVhceQaXdFZNw/PFia1Ak1Xgk
0zEb0pjOI2hel13px2FwVt4ZSk8Bdg4KB/YuIWBrmNsmiH3oX1CO8yHtXMZ8HvNb4laZng+/NjA8
qrVzjRwVW5RW7k6mNQ6P96W784Nym5INW6XwlPOnpSvWVk9HrgWdXhigI7aR3nyqAKEpOrLiVH5F
kt7lugVCstdz6XCqunaAckX90SaW3Bn4QPL3o3Dqt3ZK4yhpByFBGCqkCZ8g0kE0XWYiXrZDhNNh
0RTpgWNAAKlonP+XcdgVQqwoz3JTxEGrepWxPh4u0MABCwsxa8pa/8CNokCBh2EpYL3Jrx80sqF5
3VAdbcExr18c0CZ97st7NsYLhhWNtsmmhs5IPH7QC07GwURdqij0eOh/dqmm+sqQGMQdZjHQeHvD
ejGIGWQKkk5PbSH2GCsZU6gxZblFcZa8+A1karEINhRFBkez5xAWEIRQ4TWP7FrcQmz7xJrXTJMZ
yq2dst6YtF1phkuFWLLAGIm0cn93Ld6GOIXkZjNtTH4rHe0JEd1w1besx3fYlTVDf/AHFM7gwrXj
wvrtZM/y5qwb4jJjPT7rugwDUzGj3RH39XnI/RWsmQL6s9SdDBgxG11bCkxyZPzNbOZ0yJM82JSp
8UknaFT7I0gdulNc8BRD9M5Sj6Q9BOM8t1BOV+qlljJooSbsCTOzWkXPFJAhi8wQnpQUVZq0rYlw
9tCQM1yrQ2IqNo0A9xdq2too9IcdUEgt7lNuqLHlU+RNjJY56+CehZ7QmeE30JKwX/cEXGXNV5UP
sxxSQrGgmgHpe4cxyerSD3h+kMRCcRTV57FEpWcC6iUPojTX31M33YyUnDPbbS8iCuCSzZInbBES
ToQ1SdFl46q5mU5I2JuFW/qNjRzvjqGk27U1h5bgvUtXuvGqpcjnbgJYexdueNEyGrGZR/6lsvQR
x3nCbp6nFkNgUbdEjChunnKXOWq4/x8ycw0IMC71FJVVstXNnENi5wGsPXcwikUj15gYm4Lj+/oy
OrO7LwaXVk77pjeKmTAqmuoZM9ZkiPKdmeQRvP1SBEC/oVhzyeBSJz2mSaEEY7A/sCwyGwTOuWma
QgBvBdSLBmyzLN3Ji8jjW8XZIrOPDVhqLobOxGAg8FmhwLQV7gguuI+Hr/71you6q5Amimvu2r9Q
X4DTkXU8+9PCbvyGQcNJ5ZJS4lpxjChJpLwtIqpkPIZP6iROOhbarB4m7B0DQHJlFmBzU8TjJYva
YsFHsfsLRvyPpSE34pkl1FZA8cDJjBtdXGseId8ATve+VEl6z7SPhrvD0Y+bz8IGiZ3ALN7tTstb
n0QyBTKF9ho0va83UGe9ZpLBoh/FTGzVGzCrdaCqeZh25ZWN874v+Bd+QBtMPFdN7E0Ij9CbhEc7
vjXugcdb69EYrkzIKdZYFb4QP+CxxRW0fSmmbGodldnzYyOlr4homMcAW2/tzZb9XIsE1W24lG90
72uTff1iz/WknpAXYtXLnynq9nGgDibOVqlB14pu0mM6S9HwuI4zhIYtf5+gLqivAG+ca8GyyAjE
7+CycNOZWDu9pvuPme3gEHjnlBfmYn4RDJJkKi0RmlBicj7YxUneRxaOXNQzPmmWcE6gazYOEHNo
V1vMOoDsnZcWVLTwp86JOfR4H/lnvdrNSqO6r8a7BbKAgzeSJ7Hgk7F9Y9qwgwWvYQVuDLs+v60a
pSS+g9DfXo9qlaH4lsc++Ic0yITIrktRZJNfxOJgRkV/yrc7kjTVZvqyPF9lPjK5MuZRo1qHJvBS
XAWDSrN4TLzqG3PRQgznIsw6/WYpHbCFUinhmo/bPjWcg7MS20u+gfSgnw+FeeXHKdk51mSGJ4FY
qKpk03ba7EAONz7M9t+eHlJrFEhp357TvkK0L5ysEOtnIwOurc/uutK9PCBp7aAdXjJJcNtLCuVK
DNRyUVcqomJ2quydn4IDRN2SgOAcCtfv8l5hHJrB1X5Wn+VVG24OZ6FNtfW6rqvEzac4azyLX7kt
UeEO8GyfgPtLKQ0y8IWUhNveIkE5tvHI5A1SGYvQVnMo68BbD5C9fyuUXJzRIVhaWQf+llRFcYZJ
4u8IU4jOOUyfBi1T6tEIyUljoKPj/LQgIri5v/YZ557PsBxmFvg1G1L3EHtcgM83efa8NVAdG4tF
VEYykg1HbLZSHlkTjsBiTxipEBPaTyjLmdrlhEBM3Zt7JPH8q4o8+SMHQDrBpJ1yNItS5efMhy4R
GW2LFWvEF7PNvVEgd7I1CV8dbWrLikMedw7E1++WaluByvgp8Qs4QDnmyE4hBRARuHqMrIExxk+u
wEdVnqk1/uDm2eOBQHb/GB/o7ktrFWSOVnkwGeP241hwUzCtxgYz8XDbYg7c9xvQYZ5hF7XrcKzL
eAj5gHiGTusIibq+LwPlX1A2/+WKA1Sh5ulUsSWdAAYDvSMmKk/XCPx53Wj1NGUCbIBD88BQ88Q7
WhYW36c3+pxISAvBv1L4XBa6uenF+VeMO/EXc4/FesjgVnbSVWRHm+si/qVIH4lWgzqw7B6FUUu2
QfeoAJC1Xow90npRgnM4Bg0dAU6ouJ9UrrHkH2N2P6lmLFGW2yaLBb+zHwzZkQyDi63DU01sBZQp
lwvB6yMMNuhQzR/KjTFiOZ8rssYSh63ZYmrjK+6JaPXDechpB35tJg0C2QristkHezTxPrwA1srH
iFXvWvhGtxgpSQFjJQwsm8G6hfRuWHdSmolFWjRpGUjWB2Dc0zgyRehOUXTQP6RE8M53JkBhyOp+
LIKCRIyw8ieBjXvIOg+shcU4IyTN+97pn1Jwfo1qo9h2CDRdXk5fltXTzJVgAPZbTtmueBdvgqxA
sK2GAgXL/BODKrARczXboqgjVsm5wKnLjpe2w773UGilcwzgr5UaUVlMnjiTdikteFSr6v8Cqe4e
X/G6szTcAXmg89Ta1PjyiGTFTuT+3z/gtaTlq3Ss8eYmxpxhbIa/3TBFsQ+s7Q+R2jh5Cbrc9Ke6
E9w/hTqXQDj4enudYsWkrZEk6VlJlacci3a1u8VV2PH+/p0uq/XJgef0Ukv375j/FUDiBIQrXWff
5+eidpR6ceu5W9xOSxwOgTwsMYz2m2VoLq66XNQ4t7qRuj98hgpsTt6WSjfYFKJfyghMJGtgOkOv
Fb4fjbZhN8DOzJxnH8OzCjsW0PLyu6mV0BjelnN6p2yy6KSpwBrPcDZxY9T+2E20TjNS0Mb1RG0K
Ql79HdnP+tnEVBKgZAzkHLR++BT6FsC4N97YeIcmwzNMUsmd0ZZnp2oXUcKUx/yQoImQnDvoNWfH
QQTifwq06au3j8e0MKJwiQ4gBjv8p5Uvq+xhC1rPYFevjvi/8Erp2qVtO1JNJ6C/E3Khxspe4dJ/
pJSVySquw0uKteVfmEfF30X1Ykbek2AX711wa82BcuoXLKfcwSXccGg6YdC49spHud56MaBfg+DG
sdkaGsj8vIl3FeqhPnTZH6NajwIl6szft9PqyFHXwA0HLlE4lisqs27XWvMkN6sOokYtjgKTlaa/
N3blinbKRO+NC6atnJfjRf65GeQxQ801LycFaRRnmaJeQ5FPwX4kIpy8LXTvwt6zIPSRRqQge+UE
Q6ulPolPT5P+AhUneMPxnS6fRrKzUHAsQvHLa8DrhvuWCR6t6G+H4O4LDZMjKoeqOQ/fOo/fEUX7
ghpEgaSZJTntC9cDb0sedJuC2jbbAtxR8mdHM0hsfvZyURAnDl+lEZeLG8CmN6Eua+Kh6ZtwMc6O
9G2SmJ/NPMwb+Yn4TGKxLJ3w8WSkTnh/FxFr4zlM1/IFsKwf5EAxVQjAnsXGHBaBq9qsDEVuWMQ0
db2V6Do40mwp7HzcC7IsFzEEvFIcsQVHob0y/9h0tBGR4TvERl1cRp7adfnFlIUsDbqrGXM5dDng
lyDP92QA+vF8QStUXoULyRWjZi8PPqZSRA+aAFZOOZQ6T62PQFh9IqoBa6LN/3+StjlWz7pvIVVl
MdjSi17O5eoAK+wprlvRI0Mpq9+JPOIYkKvWsMRTkccI0Uja2ys7WHzXEXf90jUs2tOwEmjgeHOw
KIe7qGLtvB7Xq6reOw2Hz+mMRtUFsPNQCDhmV3fVj7a+/KFsl23RxUvOHwNcz9Sks6l6oTzxtB2j
OCN1YuTOVLRcE2ueEsEwHUh5AoQdO6Mt6R0DpE6rU7DIUjLntyCpGOYJGzVc4o5Ysa7KnjNG0wAP
EO8VaScBFx4QbmzFlDEJG1YSu3n80xy/2xCJ9WF7eRdaFBJRfLz9yxfcxbncM938WX5Pt5rOpzK9
/HPdLpmdJ9ke9QsZ2oHfIbwCYSUVAqy+yHQBX3z4WMMoBF9PF1oQqmrAS/WY/Xzb16AVIqruf9IO
5KmQ67B5EF8vefCX4NyJME4EopWlEAo7FngNm39RXOboR+KqxLNGYiqzP0AR/bgq2TwJShAH2fQW
7zubczbg0FQeqineeHhorTBzDYwDWkmyAThACu0ntsNhiiTHo0J7x2u82XnDr+1JChRIU0+frfrK
ePRaeYSeo3MhZqvtHmpdjcfxl1Xf1/Y/Oolu421pf8NTJSer0nm/FAB+lorruSUWW4kuajQAA1KN
oMq7PmcUjfwsChYvVnwT7iPMXb4Bqts+igHr+dHj9338ZncUlhWg4MqAx6cQk73FsXdI0KJz5NTR
TRA6sOMsoecrJ1+l80DYCz69ZNdxXC8RVuEesl0BIeZICmoOisNXS87IYyKx30Scs59oTCWlKQh6
D5iciPPB0wZRozG4U8q309WumNsSz4h3BwdeNXZzIoGozovmyRhWwHRWT2IJVg2kE3FWNTF/WhiO
4xLOyC4b2Np9O/HLXS696LtrPd0niCzm1VXWe3o3LTrFq3BajpkBKEJ2uRN7ewc2HgIlwPUiFbaw
D8yW6ERWdCJ0Wv3qwMboIMGJkzLy0bqpV94HRimc50G08CACWxczvVXG42mpVlxS/5gbF2xU6wr0
DSxPzfAR/Hb9366HafRWIejkxUFAdSO0MpipNP5aHsDt3DG9bsawZ1oM6b5szFtGahvvpEaL5KNd
qT64y2sWrUHfBBFbIinM2oFlaNViYVvm8f4Gc/VVDPGU1oOUz4D0bD3MEgsX3qJYyropVfmRpLKg
8eovOT5G4esQTCppxHHeAduqHonCcvv37pJepqMyirRdTpJ8yAx8Fi7dHt/hLrIkfPlvCwu0g9Gl
K+BAb6QZGMEdeg6TjPTlboYTFsjgwoQlNsv4WsE0ElY2I5vOw/+oAisiV3T5CBOcHHH6u9qTq/4F
8q3qBQ0mmIKkZeHPDNijn5PzGjRwq2jlGCZ+JEMb+v+HPbOgpdp5RjYemC+alPUsiy73ir7dEPmT
PFAHvDtOB4ASUUunGWM+JehIZGBziJYaqEfgmRmTE02QzNNlrjXpIgDmnvPWk6fWIY/XxvSseqeO
MjECFs5wwubQtWH0/SncpKXjGU4PZFBJW1CZxfnKAHurM/7fRa6IY1qagNiX8BQ6si5jnW16M+im
YNKFGKD6iLNRvTZfCXfNYW43MObPFedA3rBJSp1bC8aJllqJh7H8fe8aM639B12adZpAArvJqDvU
432GufQiErm1foO6c0AIwp2MPP/g/e9Wmnahsa4wgPz3NwQlkODk7vbt0va7fQ/B12lXRY7lvf9d
vRUIt61MFkU1phhnybiW7+/B3WqgeomlNyeJ1ZGyVxx9ST8+imJUoRcvjL7a4hcl28ifm1oEBNQC
pMy93/Zd+gGyGft7NOM9OcMeQ5j4wnpD/r3VCTgOMxxh9XBcpE0nsCdGjq+X4hw62yVkg6BwDgue
3aad6bCNShFt50BHIcAKtDo3zNUG7TjLHCZ7P7k6k03stW0qNhi80s/cF7eCtT+t/O06yDcQYOYH
tjSLf21tb3dS80Ks/esTEkkZugL1pHNpPn8tDy4ouMigb3UQ6hzZ+mYFt1r2xJ1xTsEQ+ZoO9JyZ
0YqYmvhtqxgCt8NUbVQIagCfryRgVxZjhfX06yVlU3qE4MsjJXeMVPlBTzfgWlzJRI+ctvFMq7FG
RZLTrS3JY/5kjiq2VuKRA6KtSXvtCcrDn7e54HY8clwHUZkXBkAuvgT5Xicz/YeLFjPWszhJp/bN
4/1ChZUgQQBc/bJJof61py/tR++tP/TBT9u4wXhtXb3u7cAaFgvAMQFOmexnhUe4Rccdz/RxYOUw
LbE2ecPD1bUEHvj9g9aVAEpFDKFckYHNAAyG42HllbqkG1jcGexZp08dbx0TzW9bn7EjJrXA65KD
nDcWdt98vXQdlkyJTu4vRH52ZaF3U30m/wjRsAC7qXh1ILa4KYcV53Ul+iyY/H7xmxNnAh1Qfu7q
0RM7NAAUZvfbePBHiSG/khJpeBk6o6VwAGZsk23Y0Wzoe2EIAGziuGssSSQnzsRw9LWX0gBhgoKm
/GkSaAwGZJ6d+EIjPlLqEfUwUXxUPF8DRFx51EQwLmZvP28fxdy7L00LvPcOMZWWAZwXvJJHRUFf
xStBJwkO5/m0RepZcIkm3PFfZz0MB0JWtABXK5FEior907d4IRsc6OeTfgPJn0AT1HmdxKot2qvz
MjN0E3k+Z6442oBVGNpgIP7/LutBk6npu3PleqxF/WCjLDH+aBCfTwBJihCXieSdsVeX2pXUCTRr
Wj+O86fbcrPsT6rBOSsbueYYwh65jB6qa9tiybx9mx60k4m1v5iBGNySRZ5//nr0n41xy8cU7BrQ
a1mqPfXY94gPVHb4piouTdcOjCXsy+lvWaHFWx1Mcj5C9EIn3IIufcdPzkX9x4VbT6mvWxJwxaQO
CSwxxtI6W7sYJalmo4JcWmUXWf3B8UACDKFyEMQHmnAScOj/aI/ks97vZJUqkLyHQEBA6n/cd7O8
2L3DkWsyNAxnxUX5oI/BWUfALobbPHlJ9CcJvpuj6p6A9L8NG0GUwUTwBUpzmAqKQpS55o5Pri82
GocavBw+ToCtl8ss5kZiqtZBWH1EU/Le/cCNn24oFqy0ZxC86FbWphjf1WDS6sG0CXX4af0x1+ZU
p3nJcesuYQmG86SzrOSYkxGWYN7yIRh18V5FZ8C4IGDZd6Yt0DKe0RiM8Ias9FQWuwxLWwemFTBu
OcLM9mr0aUp8EemIAJh6HdQH7KUq4oHSsidpBEutUw/AxrVR6SEMSebah0vYcdHCjwfwNNKkj71J
FT//tUF/4E/23G9hFri+WqkjGZ/f29I3bOmvw5RKGVKI/GCLa8VGPx6QfBJbyRutivhOrrO4zRJT
xRMlIFHRVnxgFRavvNyWKXwge6Lql2yZbH2vBSC/0qNdzeLy6rY1If/k2RHwqpDEdDtoLsoUSDIr
FA/KEP8fuywWWTRGg6l+tIMljMwn55sP4npKl8wdpi1anBBuGifpsq6/kvknqkJKPvHdT8cUvgcX
0Jr+kJgb/a5SzpvUxEzgkOI29XUsSPfcqJFJeIqiaWUvDJt8Kftdh1j9oGK5zzTg3zxEd3+5jIGf
FQT1vaqsP3suCxRk/osZ2VoD9wyWGAQL9/00MS9nZ4dO6snPcFKKB5vGBE78FJBQxSLNw1gNUANC
pkVHrOvoWS21AR2D3mp8BZIyLSG3GA6shhkoIC2SNf2SKW0aE5owouwFO4Mw5HtvwKdGTwXaFOco
ePJCHiIjeF4NW+46FlZHxalWQj1y5PmfOFazz+WIMzB2clcmSaY9yNRUYkcg1ZPYQ0KvTWf4H4K+
t4s5QqAZJM3mg9choaVa256v1y0TPoPG/dNs3SOGWTUU9jUdsWuYjVr8+XjGLqTHStargN4DO4ow
75X8AcaKvW2iLca9NF2cvxMqBV7nh5TEdHQcln1q12bGcDmKcXsri18+sGvLW0LkEKMqls97Agbv
Zd/nEgVqaA2ywjPiaMu8e9qbRQTSUbccriZ2NP7zjTbY/oQd51rnun7Sdw1stmEmgVWqema+/8+t
9Xl2k33ZKwvs9a0rq6WaxIt37YlH00olWAIp9fGjqu0iqv9v2wUMQE9ADgMTa2XJ6sd4M6tdLLkS
YB0CATFXISSeOJjesAEj9aBzSnx/1l+36ggkX7GyQ6DS0H5QvJwWaItkREPu4qlWB9LVxE9sp2ek
APrUZtxS2T+IhGkB/0sZo0VhLjKmCyrB53F7NIuhVuoz/SAfXnDzJJPv7MGnKRp7VIKwUcv/YePo
6s0j8hJGVgQO9PKIjDvhhlggxbCccSVgzN5T6Up5Jn1PFesqWmBV2bfUwZaxriF8V7WqajkaOoR+
QAmxDDYlpyBHFGSXZo2R7V0Xymj8QMIlTC8RxlFMmMjPiitxdlyiIKhwM1shemPI95Kv+tGStvz8
XUbVLN9fLWBSXB7XRBUXr9T/eCrOhk1IJe6WzH7Q4V0g/B2FBQq1FL9PbrpsMRwWNabQegSAYDNq
fIgf5xfULMGZJ45CjyIH4ihR0XJyTN5qVDLliVs/2mNkMiHXVi3VNwet7nfWoJhhuI0pGDiyDW7I
WUaHO6Y8Q2QDAW2XZrvKmiJ9FlHhmEXW60LT0HVTi7nWrzq21C1z5sHxt3AaO3tCaguhhW8Q9mPF
rYCcqdFNAGffsjOkxo0W1YfWoWo69Cqtnq1tZiVgH3b5H21okLCAkHt9Qmp1dcCobiGuQfj0LoTv
pcyYYzquLAj5+CKkbMd1QAfeDkhZrO/kARI7ugod+0gU1V4hBFc3xKC/+MfOl463ZxTaWXsJlAbl
iicasfJ1VFJ6iU00Y+cfrDZxbNzlpDP+/6jBFv5XW9u9M/haIIWwguU67QlRxTFQAAKcavNT5YVL
UmgXzFXdvMN51F1MTqWQDO6VAkN9Dn9w+/+0jpnOdMlw9h6HBwQlxrXgkp1HXGKmlubvFfZOd6FZ
IXScdNEcFHOdYy3pjuWvj1Zy0aSl6fjPi4IwS6friUTPLILUaQYsAkXfGx3UJxZHqD2U1XRcxgD3
/sAwBH/SWvUdQgzBz7vklq+VynjVAOFIq0aBuHv2/Uub+HyuZSeQeAk2TLS5hIvR9hyVXf0KdkcB
8N0fdTP5tMTojl+R/kCBQyZy1D0+uX0pNHK0wH5gGBZt4KqvpgELERFT/z9iZuUhQaOnlBr7aQ22
jhie/xNqiHxPwa4R0U2KQN/zBrvNTjOtjZz0w3JgGpE21PFr5DRdAdRRT5fjqeME9sZV1/GnFRly
iBnHvL3fcDTLOPHG8HjPOoZ5vcbX0O1Oe2er70sw9qUiz6hTDWwDS9dvDFzosD+WGUCQk62iGlPS
C9r/DM0dt1+QZbShCGFDBdRIH5SCoW19860/d9DNzaCT8/tuoMeEcj72TVwEvMLe0MfGdE16S/fq
07zAhURVikCIphUVMIoyd4EEEEGV3RjMriVLQGmaqsGpINUrkFrg5M41OYopfplC7/7qMjldNPUK
WlAPtviYBgHKNoZEUu36nzYRc9pc9wS1Ui/Pcn7OZmZHy/CyjI0iwcHJWNIX27D0QQHpuh+Irn1B
d8G9xuHQqhJY4VdTy0CmaHP3sK109MSk4rV56oWOyn7wT6UlDyFv5CVL08grZjn9eL5794xBYHN5
GgVlOhgmIyTQNnqcJzRyEOe6rHVZpMcNszSm0/TNxjYb14NrAt+yO6fzBotDUzgaCmF2edfLnZlK
ytJFQFXVkd8i56bq4YvRbPaPzQKdeT7e4KiaYlXs0+GTGn88L1M3cY2TLd0Np02/r6XXpruFLPg3
Se3V5NJCi4JdE9ZFOWvcUqTPDDgetHZO4r3lBZjgZLPqg7Dd+42+PXqrscpSXEgkMFtxievcY3er
Yv1IuZszZBGhpBaOh+ZCovl0t9L5R1/FWaG5fbTytR+9pHUhYNyB0QEMwhCDHd9L5IGlcyVkXpxk
OoSOM6WMe9eS4HZziESmgxr3VLUa0+JTWgjBsOBXxnV+Tw2tMdgBzpWFr+08/RQmAkiGnPm64ryM
3FZp39GyiFClH8eBZ7tpDrmR/iUajgOzK4DjS9lvmpnL59eALG0MvuDlZSYY46GKHaNmPOlFKRwu
1VOaqZ/DOKfj/hRUBCLXMsyI7zi4x4PPrbAornjH0VrtLGIIu0WT4FYIC/9WZgGQlh/jFK8p5Icv
gI2+xh8XWHDgxVzK1GDDEcFo+VDHwwfgAG/6LCXKp4xrY/j/hcjxaX0zB7/Fei5qGd3Z2ZxBAk0e
lxQSVALVitsIeMG5BnvbY5C+dvBraYM6pAjrCJHrOi/GWGm1/7ZMT6Pzs1BUWL8M50h09JyK3Ye6
+v5gKhIUInXMVXKPQjeMnrr2pqzYauEXLtfJtvrAcag7Kr8pzHnFbfn9Fz401D0selJkpIn4XQi2
MDBRtKHkUq8hpuXbhcqfAxPR4KeT59vTV3X2Btr1aB7azq/rvjNg0FGqpjNYKQnWWMhNZmKMqw4u
cC9eAdTUMkZrnyTiEjZiAQtQaTH6iTAZytZOeHV9ElJyLBhJ1VulMIhvmVE7IoG6j4n46Z2k90h6
MMppAgqeUKe9PijvGba1R42xI+ESZHvQ3LrtBKp3fqJoV0xlpBuhDVqNfmrEmi8umBEm7uwW8YAY
mHxqYnNoZpGEUG4L6zGBHXli3rlX4XGkPmbmHIFlJw/ZFYULunc0Fr9nHP1VWI8QniDwkB8LIDEw
4FVDxORxp1+M9lwwiiQyAd+LAA35yZsvpfllo2NX0GEzg2aoiG6m0VWbSt9Mb+2svHg2xlFUZVGR
sCKtve6OBF1BQ2kozhqyln2FWugb5odb+SveqK8bJd7se0aLysEMUnlWg62LGuEfl3/WnAGftVH6
zPnWrBIClvlseigXFgUlslMDRChm7wkxH6PyRp0nSumdKX7kjiaVp0KxzwHIZ2F3C/cFW2YHrxfl
rkltfG99My6I114zpcnN5vfCEJaYd3vrGkLHGXIL4TtpkW9TSjTVz59/1oc7r4ms1fC7OayOpLgz
TRUw+RdhFGMLBMex8LaME5NeH1n9Xct5S2PaXbQu5UNzAUE3FCWmCDrmICb2vHcSRM1mow8Xtkkn
EdsGSpdXrEwgbjwSEaqMgozCtQd5C+YPAdXaPub8GExJwUwWrbPgxcppSq8ZqW3N7Brpq62Xns5W
EwGQG7kQE79Pry+GrS4YQMUi5+CKcL4m6cIMJKvyLYC615QsokFX+wd4QmzjTuEYiAPbMC7Z5aNy
NBFO0jmCx60iZsRMcXqrp7SEzwsSQ1lRZwBraFzLBhaxmIp0X7ym5oMm26vmIRCrwHevlWm6ikja
JO58ah0rqRPURoFWSJEc9GInj9udQAAyQ/mRgqRONCA5pi6zARPPzKu2SuGLFyKtZzmlGPtTWObf
ioOGHbv+aAXHp1bSZgThkioIgbj7t4dRNBsYf5PIK9oa9rFHv7OB36uauaH0EWFyMoZnxXiqDBjD
dBXarsOwKb+o4o2GpQgDWvznH3z4huYtiu3qOJ5FB1/KF+ItOyi51IcEb/AiUjJoTIuQs+6wyBMD
yZMYmik624PSqwMu2MfmQZM4mZW2esBJsfd6wgR4YbVQKVmQNm1OJmYYrbr/MtQzM7JdsGDwIjmL
zwF6Rx3EcC1fMsH77ECAOaZ3hLc5HjVBC5PTHWM+frMBhRJszwDYXwaI7qDg5tVMbZaYqGxSzwJe
nyiP3P/qkRKsHEyBehIKM0UsucZ2fSqybHeZXiBZrl0HxgUOHt7gVbF2+b0Uc7wlag9fmFJ3xKoN
neFvaL89nTUPnndZkhKnOzuZmW0KVN9pOiB2iQq7r1lohTAEtxZMD2Icllm1uciP1w/IdoqcfyXz
eKq5yaeV919kdNdRDveccK679gXILKYuDxq2EpbFB1Z0UGqAkMKGlgPX/82ds2UGlf9Zj1TAo7DW
rDra7S1NMB7a32zFHFg8P0/pg5cJY4INhhBzfWQp+1oCkwvLjAQ7gEUFnYv1W4LOrvyhiMP1+DJ9
OzF+ggBtsjoC7chIYIu11fhBZI6f2H10Zuzp13oT5gmymmSFBoi9dWybr7u5BimkFF+I85LbGfly
gQDiAm4PQt3zlaUWY9O7bKWH0jBNkQ3q2e7cv4JCnc3eok3wlxG3XYMjZ2ZgPKPFda0NLcq9abnn
27QEyw1bCRIlGj5lV9vQZ+3C/jrshTZmmAhTUcvL9f0Xe6SNeRFNs6Rruq6o7Pq/03Pe1qsbGf56
mJ2HPoMaS1mZf9JHPY0MV3tUGx+lyku3TIw+XFhq/o2mhavAj8JElZlL01xG8P+uOz5xPBKmQfSQ
laz7LTomcDbU8BEeTj7ZsKLH2lLdBB1p9kJ166WDnCwaBYtPHfbHlQ3R8DobHCL4ST9HXJKVozIt
Rfxh1/5JS/6KU+asbyTNXfWjuTKZqgVHJy3T9NMvRS/LpK4UQ/c+WLjS42ZOtgCKNX2rm+m6xcWh
/yKwzTHAVNMo0MlXL5wxwppg2BOisf1OdOETn9LD9ZKloMex20c4b/xR/e+a8PdhBQ/ehbIIXPi3
UdI/xNjFMjlD3j8LvMTp+hgmtXMPKEUZQYQ4y9gI443d19K5OxxPKXmy94OywH0ZpynK2Bp9TtIM
q2rjsNz/kMKF2smG022DR6ACrPDM4pRTJDmAjE6gpwS2bBYqhzim3XCajJb+olU+9u5rt++Sv1eZ
x1O4CNAg7zoCbuS3I0DXEgqjjpVatZhEwpoz2GzHM8WCeGzoDhaVQqxYcZ4e3pXpBea6xw5rK6q5
rlLJOJjre9IStS4MMZnylMsPv1pUR+WDBnpQAn35vYsbwUq1F4zHYUzCc9o+/MTfLkkQWzEnU1ED
IPXN8R0NvKX+l/zsSlkzxTmPmc4IPoZ44MiN8GxwOlu+9s3qVKruBULZtKqDRiKPTvtugkBxVTqv
3hRwMtsnRIz6opfn2iLL9OlnBtuNfcsBwKVtEykqMbxlGlL9c8lAn80JCNpODmDG+u4XCdPomI2w
umops0VMVJaLIuvMu9LUS7EwrzyZ/j5rpUqXSpNY8bm/M5OFgBCNwEFwlR4tIVapCfeIe7AYCiZV
88Aku7e1Gt+UlsVc9u5gHQzCHoaa+ABWrjkNFHwvVeB31COo6FsUhlMpU32yry+zes0wndmCFmUh
DtFR390njV10amRZC3xrdHB/S1+HYnH+y8LZ3qBpiTUY9svsttkG32beVVN9pMj7nPw7eCuI3hMy
u3WWt8lB5D47zBi12Tmdk6KPju5hGVs34bj8qmplglPSZ+29hI/9UwnQFIe5hSH/ynUWz2RCnPyS
1UmEpERaFsaN39Bj50kpIAHlF6b/HTgUyCGfLgG9wgquFqik1lu6WMTQrsBvtSAbNavNh+8JlaLs
DH2E5WAZacN0DT5n17kFN63K92EmIBQo24EvSdfnkY75Rw+2Q35Xh9vM8Ryog9r/zylXiJkuvOHc
rp84VKmGi0xkxy0/CB+13hYZ1/PWOiB1Ztpsg9/0OGCnr2b99dPqWJs+p7Bhdk9HLzGZuy7QzgpK
bw/wWmsqupG7z+qefydov7h/BDGmUzA2e07sUHwLEldKYoCz2/23Phap8Lvk3zcLHbvc/oa6lTAy
BfNg1wO/wB1+yTZ6PamCPrS4X+xnTEtb/dSXTchkPgIW/H/n2K9YXpfvsIwKXY4iQ6r1wrYbVRmS
xL1uWfAxIg6vFc4Eaq5qh8kJLHLo8ZaXoN2qEJml/7EGK22MPPsvEpHYLdUcaojtppd/lFl8nmRW
sc8XoWf/5Kaxnfhy/vdreAfeKW0BY40JQTOaOBGkvHdv7XFiqstC12JvKGQomBcQ03vjK8BdW/5Z
FRV65hpE7kljw4vPP+fxfCvWInq79wMFyZjp7+ZHwK9s1qbZhx9XaeAxLd4/NxQqiZ2j5xWnt5ds
0iw/XhqgvNpPqn6NdaqzyNbUuF9wr+/6M8pcmE6Tz3Kr75z+3eOvOAWKNJ330DLZ9zkMTV7nCIYe
gWUbDgr1dMaoTw3ONoMQqyGyS2RD/WfEfLcoQ7fbffamoVqyMMgm1cz2rjXJ+x1+vQNKRo/JAeJ6
o7f74/jsD3kGJA55RLxJZ4veRG/Rsxht7h7XHrRtxGlv/FRQQQfmV+QBtFRin/V+5B+LqfuqTWG4
n+iak/+etY+dEZl5c7Ozqh4js/2WGnMKz9eqMiUV2TXLhcVIKu6n6ndNe26O9gycaxyaHafdNtx8
NB7T6elA2UYYpgAJvVUMiDINjjydzcl1fhDlJIu17nNZO+aB+qolpd19nyF7WOpMxAzvxBeSwoHN
Br8V2aCWa/HpNol/wK+vBNy9Pvgl36dHWBLqwg6YZfnrGa7jK7E8tGm6dMsYkePAUpj7i0sOSISF
gIDPqX3PkzHcSK1DmPNpTnxOMjsciSwV0JG56LPFFh5Obl4zmsOXW1fbRRV2eq5++36Ac9TOK9Fx
YcAZWU4Jj/Ktghnap+cmLMl2QQItbOHYpWkQCGxAVXmd9VaqUAGs7twMWe99wpMmQ1auvyXG3X4g
K2Ir0UmZNvMUivMkrC2rcie7kwkGEsQhqo3H4e3/Ai+V3tM17TYmlG5E4P0xdhJnmROb9krUddPJ
Djy5o1X4Ja8aLSlNJFNUSWYbpr0argYPzXG3N6gr9pGJj64tN8Au6Zr5BJfiLntd+7w2k3tqPerE
+CXxE0aV6EE4exC3tT3NGPlrH88XLDUV+V10qiY90YBXcSQt9j9e1diSwBpAfvZWqnROPWHcsjAt
IkBgXcU+oJ97zpnNHRu2JNMCgQfy2VkLRyqN/sjl54q7P1j+vjyz6G8RcvUlyKOBVpby9QzhXhil
mCPpXYAs14gxfagwADQGGg6JvJT+24Iuag0nvVzglEQRv+rvS0x80o1l67IqqNlVLfrVRitNJQiT
YqXT9PnTTi+gACddCs6IggESIg1ExWwzNZeCNGiormLY9NIHX64N1NEUEwfRaP4fFja3xNgasd7c
IQV/Fm9vL5tLAta3GFN2zC+bdwWRWeOAgVQsCJRTS8N0wL6ON2cuKWFQs2sm9UUvT5bmpSrbSBX5
s18bser/ysJnV1ZaP9An6QicElazBvhXsJ6RR9bvVZXCN7pBqvM031WQ2KxEANRq8EG8pEZTI+M9
zIDlujcgU5vex4n+e12OzLTFMF9yK/CQtdyOEkgC5zUyP5xqk20Jyj8XCHkICHGsqu+C6qfw2BDf
YdEKf4aOkobIzKmhUQsJltOFRhhuP7u9Rxow4yEcdYvyAgpji0f69O0nT1YGp4zGOy7NVfiorjkb
efi18ezQ050Anjyv3BDJNhnjF6zdVAEZLybfv9Gpno4b3WkWJPZh3YlZegjfqfcc5dZJhyT+YL73
ym3FA+yUVscFtUK8bJIyDRHLoICXBx/RTg501jSepDBNq0LhYeFwS1CYsNj89BLW+Sm26oDfEYOY
hffvzD/ql+d3AZ4uebVjVaU+uYl1p7VWrw9Jw8VMcI80Y6SCUQ3ip9PyLh+cP/pFhLaXau2+Tjd6
4NtgttPNvasT06kd2Gn3Ytah3n8cAXR/55YUBS5gYpNzq2CpWLAQON7yfs3BWlnYQynuyp4Khh3U
zuxy7W2Ay9x1lFRZ8NnLjR6x89FDLQZ7SN+xI3wlDZcbD0/JjZehfqItNKhfaxPOm/7tcKYWMI/b
/qRoNSLL5t9+d3uBzInIuLN4gfWpx+/87HvHEYIzmDMN56nXPzmXRsTF9tMWct7dLu9kolHSkUlC
NBbhp1hNpaw1jK8q/weWUjOCk/HRaf3J7DJVv2NiwJFIcLbCISBY8zKGTthj2y5k+4sFXpldZdcI
PdPKrd+zMMChqU+bZwvvqrT8KMX/XNTeRDF+fdFXnwA5aMdyjp1Nz2s1KJHdg1iQHNzhXMna3ld3
sL3D1G3nWMBDNLz3xTY5q63rO6cXC39D/+I7qgJ2TsLaNdpHhjny6AbH3MscXJqjZUQpijsMFHUZ
3IzR0zqCSfDB5pGjS2mjOV5USfhdeWRdGHypCvJ0s6czp9qVw2uP9NUdqwO5mLtlX3VPHacO0IL7
KD80EJO0luHW+lAIIkumlAIT+1VcU7nuUbJPyRBZPS2ApoIeNBQWVoW3jcrEx6vxPV5Nd+RC1FZY
qYjzc9192wUhQUmu7gjaKz9hwwG97VDJo3WDAu/MOLBADtifYM0f+SZ9FAfZKVyOE8x5Oe2eks4J
iclNrU2QBMgWJj0s9wNq2csX5LNir6pvhKKYFxj1ZwZr7kWJh+lLyIM2m1lQtay54ByeTQa32tr7
62i3+2Swjzz/kegcQKWRjWy7DEeh/M6lY4NogyXrW6yvfJEf3Lp++OPSF7qsqwh/EsZSmwOAL/8S
U4zGNKTDK5DXjeFkKwZR9jPw15JCTVpkTPP95l9f2uMFNW32e+/Bl/DXDRouUji7JvpAGFaaysuc
ezfZWBASfXF9sNw/EmSpfUBI7z7Ra82CAiqfGemIXrvCNOZz2V4u41qamMTMutBuAYQ2g6sHPBN0
3wlolTLLCslAYZ+AWqjZLK74pY/ZRr/aguF5Uf2BC6uHH59LKRNJdHaYoYMKCo6FMux0tK6XyhMp
kGl/c3UTATqcTfPBL4xtNtqPppbVuLHAtwDiBW5P4D3ZVvFdaw+BrLdX71lPii2F7n36I1HtRb2K
ECD6ELX6NF6Vaib2D0Wf4V81qExFD4KkyGN1mJbVmud0JxszYGha5jxjZS4XZQM1+vWAmO4xxLSL
kK8LYi/i6ojA1nh/EcbpV0Pi9JtrV2u4O+WG1xkQ5t33QPDwzVb5YHJBBQ6ac5nXMoNSKlpTmR1a
Uu55ELLjwvig69kxBC7RL4/7IL5GgGpdAxYfy5CzjPtVFjyGFzDA+Tu/tjEtna6ANyqKlOEYerIR
aJTF8c+y/uZR7JvDjVPPD1Xt3lbF07a6Tax4IMPBFUYCTRgVGYTjwZJ4HIXDqHomcB831j2QvgMu
cM5wR6f1v1iuHGz6xy3tVee84Ipn9fxvCEe+a/2Dxb8RNDtoUazBTN5O3PJ18Eu+CYC2ipKWKZ5d
4AAVqXEQ8a9vsIJGZijIyEo8thf4yxd1FrpSH5yUcZf8zdxpzbhX1sR/C62sctH/mxv/sYmPMQtQ
vvBxaQmp07y3RNdXJLzK3UABfK4mfGi8xghTyU+5uHVrepKq7UGdvWSsFGLPeiEYcCK5DtIRLUAE
i0gmIbFtTILb0aVzGOUqqvcqwKW7HHpzKpM94shTwSrCvwA/3UnfccLiKu5CACkv5+ME2UYnRuzn
BNB1kEzraQ8hyChY9ajLJFVQXuyXaCqb4xSvHkDFUedcJN4BtsUD0iG78B5T8Mz9S3xBDGxQ/yC+
oULyN7aovmI27gaWFudmZOT0n4X0Ks2g6hPYzswusgmtW9CAF5dQAA8j/wbSGmA/J+hRl+iZu0LV
0rLouc8HlNnXEug7kLOmslKkDKkThVdbmMp5Zl7pN4Ps7bdf+koMhnhIxqhAnLaagsk/1Xgev9AW
5tFK+VtBZ+93hTFrqjfCF583U6hLxH3nbR4hzwsQDkNxud2yNaVz16SemrXXJeeAa3feKayTn1EB
zv51YKpGSaIO74T1Ug3dVlH3LVAOmI4DzFTk4BPuLMF9gpovJpt/RteqE3UThSz1g9xVyKHSDtnM
hbrtWvkJE0YLJnGMoAqYzExwxDdP8akNqBl//SLU6PzWqghTvN90GL2+UejOZdzUdA0PjIkNMY+m
DiyT4jLWklvskwM72bRMyoJEH7WwwOiyGTLpO8OmykPgYvOEPUq15ZgKak38wn4kS3JGhpGpjBvg
zbTfO97F8rctDEtBvZfDuxe8Tujsc4k1uAL7MjfFSE4X7/v1UJwRh+JglPKrtq/5VbIVYX9A/zdT
2b1nHgw75+ArIthnT5s7xOJYiVVPUvtMMNhcDio25RaSXnN+DW52lB8ulLMDLtA77PN/Rm6wLB3t
b98au0NyZHQ4Zgkon0eTFscAqOZFvfxeWPKNr5UTFWXCpqEN9zuJ9rFH+szBJK6esLauxrwiSOMY
BCTEDghsl1Wt1vHOLLF28X+KyMgEHp4y6kjqlO9PNCmCbZ1AO0h/k1WWo9VD7trzp5PWUKWZw7yL
Uv1ujt60SjE3J0eBtAwW19h7vnMzrBKTT5cd6gRqk1MKfasHTIhmP9u06QUQAwibpW+AwPkef/7S
JPxiIIpNWpnMdmA3qT1fGJGISdp/2LRQzO8As3GxdCRdbghY5/3164KozxgEHAFyHJFY2Gtm3h1w
oNox3AcZ3WYlqK5Dua1k6UpXSxpmocEnVcU8cvTfzmxSGW5lTOSGQen518i2fPNMoitVVWY+jp32
3myYskjykDVviffgxThlOTP4wzj4NLCBYBfHl8ywghhaGzzlAIM/uc+kHitTzEmkm9st11CyDd6w
Wb+Vkc0BVbLKF8tUmUKYgcuP9LkounU4/YaH/z6d/GfAM3YzDhq8W4XhHRLRlk+Q9Z129VU3hP7L
rfxcSyiiZD+7zbdsUVSvfboGTIiLZee/rfF5i5/mqsfJkM83r8Huxtc7z3roT5YWO5CMd4N4qF2n
lmO+ooLF6kbCYuzjTf0CqUJCnvmUiGHvGD5pyKObttovIEv4+Pmi6xsnAWwpfbEQGL6aUrd5FX6c
CL8pGaxcQO/7fQIDewcpQVJpcJby+XnBU9sOnYDrFwZpLXjgVlC1ZzcYRbZEW91z4sTUw+ZCtwGi
GZWNq/q5/v9xGtPdhMxobuZZngbMUG9T9qLyxqjolPn+onK8c5y8J+W0xyhzH96dpbD5F++82jcr
AjdtLLBVrNzAB1cx9zI9nxbN9b7WeJPNd5R1QOiGzGWihTK8N+E08l3rZmsoCNIltm8eLPPjnHj/
ueSnxdtrChmDoRmFcdAx8PoI/6kgAEZg2k6KKanjEEC83b76wQ7AmdcwaNiVroOVVfC6VsO7KTfq
03KaX8d+TfYCuRzxJp0RXFHR4e4YYAmpTM0TAx+EtzFXgN1MFqiIfsrxTku4uuEOX7XjhXTeWuLO
Y81eU1IcDFcFw0Z2LQRG1q7rCGRuGnRmyvcB6weGQ9TzvKED3wvbDCtisyc1zFTfB5VCqPMgVou2
trdhn6W2WsebIKFZxQF2WNA7AxqNlJiHiVWqg9aY50/2eKm9r3fa0A3Mv6jRQLYIQNqZweyVrL1C
oa1+vVS+yW9srXEr75SAcyXPDGX/xOXDsVy4oOpVVKW0hsRrPq+dpf0ZIUzqetelZ9kYOFZkO7O3
uEedQnYv6vjc+G4JPj42MybCpeFbV6FJpJxN/sSW7SxritNY1t/4idKg2BlspCcvz/gmhUyspGBh
f8xn5WuMLkMY+DM9XzyMP8FMsmmjDkkuMMK7XRh9zHVrLO5ClTCac+SidrEofJI40pYXtGdN7SeH
LJwdQeyM+xUm+ucrbFKjl5TgsEe76SH3LrgNWXTNPesL2RHEbZVWTxKHBAT5/P5rSsA5pe7sFSow
k8xRwRo5cJg8q//k1yMUxXgd9DikopjmSqNTv3IAQBEsKKS+v+ehG4WCaeETajdV1lFj75HjUmBm
uU/jjKmIKpPGReQZkNQeBn5y30+0i3WjjMb2RHSHXK67fil13isSJfWHSrfAIdm/2ln9ksiEEtEN
Mw/mdffWxfIJxdFAEdOsKgK/8e1nI51q+jjQd+DfNZmz53t6gZXsIKESUrzfTiTaOeJ+V0vYdVy3
swCeNMb4xa6F9brFD5b1TQ6Nt6KowUcFaXk/f+K0+bAsGfeDAdfUaZqZp60Ae8qnV5QMA59p3Y3+
M2MYWrZFn/l5Hc9ayZcDW5E9PjmdpVB1iBKiyTKBMg/inB6j60B2wfxCl6ux6UV3eVDmhec2syNi
IdC1uIJJuNVwl2/pFfsyVpP6jIoxPVWRRaMAxepGBJOkwQVQzFuOOOXeILbzliYFEjJfNXiPgv+/
eh1F/mAkVZ8FNT9wOFQtVfAeExNtlctHx1TMVs7K3dTiF/j0jtEq0cZ/VnutmMzRxtno63x9PyM0
uWyopRj+dAzX1vYh9D85Bvu+bJQKcOSTh5acq/RHMYX2f63JVp2j/BlqNfWIimIqqbeHj7FFPq6Y
ih+Qbk5yFD8jUQmCp9Nl2UGyIyuRwc4O6jiLSjDF6hvY9VQufRoIuZDdaMNFCtNMy6tW3n7L1lEA
YRWmbbvzYD1szvZdHjT5zlMc3jBfswgTwZ9h28NKSvshvyLVQ69GBXoKLLxMUPrQymGGdzWJQulT
v6gQgM41l7KH/EGNbBWIr/12QIrOo2uIUkSn1p+Wc5ntshouGvgOndmDynSbCDGrffPe2r3vMoio
azB0PzUqnITSoLa9jlclH6NxcyM7cF8kQhrqLcVEKSuyf7PO23BM/SbJllBBXkR2w+sM+XzI1xjG
KUHVBG2gK4CnXkS8gHnErausyfJBRbgYbsjNchpbq7+JG1znSoohw6SYqAEVsQeYvcOUnkSsj594
IP43EWbkWS3Cc2Dp/e6n3HcFnSU3hecKgdM5jpRUdTSEZkgMHI+aA4cMXmeVsJozHE2BP8KE27kH
uBLCsPkHBRYWAwLcSwa525sAil+kL7GLh11HLzYskU9cICk/hwvCCuRUe1hdI7lJd9l4oLU1Q4ZB
D20rT1l/ZOwU0L/KnlQs64K4BkqEY7rZ2XopUpa6C93bGO7vGFPFYH2JkhQAgQMpPtsC1lL6loth
k/Uoet8EVOUG82/DQ8mcbmzuMWQYJ9CxgqUHmCdx+nTwsUpDYwVdJhvbRQBkk3c1xod/vQ9AmQv2
YFPFZ8NQJLnoBFW75PPBZ78PV0NR2l9mvA/wU1c4h5XzBGFlKYD/osWSZKcqe4fXh0nijlRhjEAm
zh8xMp68+26Ki50HZFdJJYurf4ECzbJHW5bQO/TES6FIoiD/da684VcpcTgOoA1U5DDyBBCUOAz9
DP+I+7g/1wmM1ts3GQXTv9eMLhqKAy+HLozGpYmP7RxFZ4XnAMhh60iirbSoTmAjiInyPwIIvcGz
/ZAKzWEdU3BV+jnmt1645YAW84Aa7NUYihDgptBCcYWX5PAajXDGdC9O9b9u2U8AcFfKa+ruiAiQ
T2ewlfRiOCJ8T3vW3ZvnRziApKb28MazBbtosUyxFphcTKN4g1lSbpa6SsMOO4wk9E1R+iqYW40o
HeQ5zK0sq/sGsx3nBD2W+OjEWE61rIwtor8St4Oa5GoqIKo6fIJs2m4C+jP15aG7vT8TNQEhfDDy
l+F9vriKkhx37saarsLvi1SemtDD/vjRjPB4mlsSLAVjO7YMBN21iokPeOc0JBQMD3jKfMR+g8P8
GwEv4t6id/UV0aC1kM3upy0bzhJXAP06KT08hJUIHnLbjbfvQa1bqn7uUlSrT+jvKNcTiIen85+p
nW3deAFj+k9iWgqJW+5nd9KPYSLU6fh+2TCWdhO4+F5zJfG2YVXf2V6et5X3AUPBk18rPXFhXD0v
vpiFsIyQ6xzNUyuygM0qG3EXdMpW/Gv6L2RRRqEZHJKBdurdwY6jBmduMXt7017VYZ7h1fprLmBS
LiMO/aa6IxV7GtSSdAPyCNgKgdhxwn9cbJsxePpLflmCr2ni1nBa8Ycpkt+7Cr7H8TWdQcndX1XR
gSwLYoo+rwTcmtB2KgMKtSCSNsOytyS62emIcPi/3xrPd3Hfr4BjfRhhKWm5jdfD9A6YXGZ4cG2H
D1sPXTje/Vx5YZzV67awGBk1QPX+J2bGSI478CjEZdl9MijDcmJkv7NBD4fPjfzsq7Pt65UJHdB/
Mdtw5tluq7DgUB+yYZ7j0ptNiuf4uwvmU/QCY80JugcbaynkG0uwizQaRQ1GGJfP4bR7saZWeHDb
wDU9fWjGDXK8Cm3/Im762eyPcjf7/f609Px9gKGazbeIDxna7EP8eJ+q0AuT7idZi+7B7J12g2Tn
neNoUvvOCzNhm+i7q+t/5N663gpdpG0sSQebIJqSow9CeEB889dAPjv44G8Mmcfww6PkCgM2MLQ2
OUofZNAaOFwIurCV44KkiM+Wfm+s1btgrwq+YRiLbjVVaCRp5mRIbFw6MExQ+jJ4lL15kB+wW8Yd
qcUrqAlg5RURat2HaE2Xvf65P8U3smm2edI7hgizRHKynDRM6sv5AVSvMEMC5HWwWqVxeV/9Ajvv
Y83zVaioxiBFYBHJXiIVjCq/1wbujpy8lwrKsU1/CHzQ4WHDibPfPPe55Uke+eAMHYXcyxLmYE7N
wsZdnKNL4NT0bVZcoZ+PX3oKM+S9qkPdFiwj9mVoOgzcI5fAl2zPyP361rB+3wEdox9Mxqp5lAd/
4nrT2neOWWKDF3WxUPgXrukgF0bnuM6VRsM4oPFhgTi5QFIKkHlI2AdUo65ijWrMzLsC4qCUV2mU
JlZG5e/85+6fkNDKrRTwfpNtSb/WI7SWplVsPtHINdl5bfF6hxP9QkU5ERj1R6T7OEV6csw776FM
bctEMi4IWGSVEB3m6ruZSfTIzXVIS3LPRZBCsTNtC3ng4wwUnw7z2AiazWnSx2/Z0EBIwmAYn13u
FV0+QvdVsoaIpIXxzHbLoJ//y5R5fUd4IZqO5RZPqe5yFA870aES0zLbR1jK8raOw6xtdz67TCLR
G1jBJhgp6q3xcgGcT6cWefb8higzS6GhvLYwqIyqD44ppQISuHt9i02R8WHIyN8p8NrqtH3XI3cQ
868rm/kgBfCibkS+3GcMnzkbJvYHItdwVAM6Tvwyvw892GYreQTg79NviTbbM4KZNXlAIstVH5BA
5DPTv2a4XxFMqmJmkXGomfPpTjoFeU1Ewj7S+Rzvl0PoC61YXJwaDFVloBmA3zyekfYtYS8tB9ZZ
VaoOIzBVNm9mGZMH9xo2eBl7BrUBdVtKh3fePU/l+2MU5ODHdHsZ9uwbAM7q2tBcwMJDCEG6+ttS
nMExbnmyOswH3qXu7kH+Q3PNzlX2nGvWD04+ybSsVcV9+kDEquFzXdoTL4Oxw8/GymS+xUBx0HBa
jmBaPsMoooc8ml3fn6zofWD94g0Ra2AyC2/lLaD/ueQCmg3XCZebzngbSYq39VIDFO0gBRse4EG/
nZRvDTJ1bf2Q5HA9cUPNmg8s2P34Vze+C2nzBgbe6orWRYByDancaVpbtFfcWX9XIP2FVIqzXJ9z
659UrhshX899AQG5MLjxmUAABykffwjvGGdyMkLMPCHof4EQXXSSaF5szji/wKps6KUp6y4slo0L
73/kFlUp1Luy7CLjHmKO8HY3gLVGd1lwXp5aN7NSAItkSrdQe+ku9u/+YYC6tkHcVSEl+a2mvl1J
A1aKK0LBOCnkBHytYTY0/k+ZRbjTlUzb1M15TiOtRZbnB+8+AwONbfiPnNl+kObJcwkeLvmSAKco
HQoyQYwy1yyeGCPxdfbr8lw5IwKrLjFhrbDVFxfRhdHWayZ0YCAWeB0OqUWEtRgTbX74t6OzwlGU
sIshGyQjZuUKY3t7QH7GVCQCihqjywj/eZeGktbXoq1IIA60NrphRzMyFxL+QvC2l7ee3fRtZ5QM
aHUlPSQdqrSzjP5/qYe4sLkemYA6qRG9CbvDhbC67mHd7FLJZHBT9Qor+aORa07pmHaEGxcFusuO
mqlgM25Vat1TFUNsYbxYWrd2WcGsMskYd3xMHMxHu4VZ3Fw518MXq/JItTocexHvlbVu4Dfhz6LX
qbhq5WRio/eaNpr4KHCDaA1FUdGMkfJZUSMO919gZK/MUoQ3tCexwWiwQavZEqeacqxrg8uebRf3
YzSw9Hdvju3B5QpODevRflWcD6Xg2HRjnQDJEcOSr4Rb82G9910KFY5Lxe7GHhQC0PORO2JpJQRx
pvH1E9cz+ihN4kzx8jQcubL0trmolnywxMSrBcrEMPkWSUzF79hva92n1lJEOBpLOxlcV/xZqfCw
oMBmzUdYp9IH59PMWIC00O3CryXAEw7vjdsLsGjaFOanlRDt14zsRdoAv7FN0JdDIf7WPr5202Iv
D8gGJplM2OVaM7jlg63DuTnkrx5c86IUsrggMKByDuNhNbE68iuTaOSh1Y39SrFlOroiRpd7Mh3u
CNPA9OdRZAKK/D8noYawGrpi06CAMYlqhLd1FMpRgVgg/gwIW9BN7422+7UoORHg+rNYIRfh5eV0
YTvZ1FEWXsOZ2naBlAWILvBILwRCrFrG1aQWgO7QwOSoTGU/u+J7bMzHnl69ePx4Kilp/jiyThTo
JPCkl+4vnhEEZ54MMbUY9ShfrQtaZ2+3c9Uh4gDA93pQE6Z12DU7XYARJdBoqN+QFAMyFeTRUY8g
bDkGcf2LbSJiDmNptDembWvc49rB4ZyxXvxmfm8O34vBgopA3/8TsRs7gqd0vwqt9znVJsUjnbuV
pDmUVgD48JkC7QfRYiRetprLQa1YWicsVsCkaw8MooRNc/Ri83sJ3hxqj6fgNF6ppp98Uo1wMcgQ
JdHTj9fgeJnykOeRqC3fJL6qkDFjqbP+p9S+LJrpc0xbkKBB4GtGOdGL4upcGU+7ttksjr2nRIoi
QSyppwOS7KrgkesmQ4qzgKeqp2SXswRfCJmiFnzwmNnjjdPnFveL5x5I6S4kVd3wUIroojrA4Yyv
p7n7nnYn9nSuPWOCgRkgauIAe6CPOcBZEkFHI8YYzP2cmgHHKaUkC3LJ/rShmYclAdU5vwTkWgQD
yk5YBYVJ7yqtwQk+2Hti0sjpV2nlJkfLmwSGtscvXbdQKTkBAxpiyPhaJOQqOI007FhY3KJkhQLm
/RTBsvJtRFKuXghZsdZFseiVsuk+ZkLrrVEi0+ckmWh3kZXB6+8XQXI5yh90164J058uM43Gkt43
cw5VQnIRqUU+81JmZmMy9qN8zvzrJC2AkWlXdS6+iBV0gcC95fuF4Y/5pm5RivJJOYGT4fReu6lU
+tyvrpXFUESHmPSmvMMIguTZqHFo1cjpi8nDnAUSKAldCK6wYAJ5ICh6ertBuIA2SpDB9MTBl9vw
x1aisctXKyYUUL5JLFiRg9du3OcwnZemXIwpH5WePt6stoaHttZSpR72P7JoFA8QSs9sh2hPQ7qW
c8+qZn9iWU10SGea4II4CSvifIjtuYD01+PV45FU84CSFgbLvUbpE/ZtRYfQHaVMY8ZvLxN+xapv
UcTFa7LjgT2MALPLC/kI8Rlb1KxZP7TjIwC+pcqg/bEOJfW2Fn7+N0MMhiBDNcji4+X5bJF4vzY/
GBEbj2RUHBJD9cR30vxJh+kE5YMcKUgRKRYrxgAYnE1DmehEgbfSc7p9iZ8Zkx835QurWXaQjEhS
GhVhcpUPON6cFuMXfxo/SglxG72qB05yCaUOj3/NeoRx+oE/dhcntpiHIubl14pwNyXuftMkuuQh
hN9xQ0fjFe3IdRr29aXlq3a5iajarfoISB4Acc9U7tIqDRkHG1iJk+tI/QNf5t8LnohzRTUqtxRQ
3SoSzCyiag6VPKOxQ84ibMkyuDjA8qsDh5IR6PU957xhBKkzx2oB1Uh4jIw13UrBpiW+77UfH0ld
yFA8S2Gr0Bfs3eFxr1gEcUY5xswy8pnqbtLmoUEXz8F4RtR9uAApLqlivvrylqzFCfdrNKWU7Z4C
cHcSx1LCmoV7okpFgfsy/2+IbIq+OPYnGikAbSN034lQgp+yerQQ/SFS6w3AAuvkbK67BPBqG/rd
mQim5GZzd3aolHJu7keyU6Bf1VEZB9Hbbkx1i1Si1fWQaQbE9SizNYHOKKouYEQ8QhyhkqLQ4cnC
m1klDaETyko+pdE+OOLUDLDgG2WkkR3XHnQVEtEAr45iTjY7ev9qOLQWwYYAakuKX+HLum/es6c1
W6jdfx7/C2q12vUIkW+D4amYZ2jujE3xgsg0eXoiN3MBQ2ZM20BCFZmJ/HXUdnraPPXRgJnhWHKQ
Vq9kd7hj8gc8d0nHOc9R6Q9sx1vVqu+/14KMkbWtS8nrIgNWDdRkNsjEFyG2zlTrMhWMxX67z8RE
rCsk87oXasWCaCSQN55desRBMjrFIC6AnRqzQ0gWJfSxNclHdUMWjOqVbfaTbpwsBbjBYbOa1zJw
vgLYjvppNMXzYssf7La3tkx1hzixDLVEOwt9RqajBUU5Sc0Thw12J3RbAvtvANBI/R23ebizOgNM
azJ+5V3XCkfp4yW3vNamFy5pq/SLWhkwWZPF/Sz/Q15lgKJZf/uRZ8BR2xo5SuRR7eJ05o7JTSXF
cY4CvVylcOq4Y62bgxLhhr460j5ZJLMJLRYLxma80uJZ3dDLhDdL9ltLu2N9w+yYqWv5Hu80LYi9
hBq24vzKcWwp+iiZtPAu3Tx6WeS1Fs5Q1F0gmL59auouXEIn7jn4MPrtCOVcko+EqB2V2bCG+QIR
2hz7hPWMjyPdj1GwNW0gPXn2j7vbB3N6lk3bHhQbF7rllqnybFiQ7pNH+iJ6pKDQzCcZ525me6XC
Krwlnb0gO1qgpAJcvUcbmbRg4R6yqYpCZ7bweBsOjpEEI2pwH3D+jb7c9F84NXjkKXhWtrabdiBc
lhzrDf/cGevn+l1Oaq7IEe1sZqQkEWzpXj++5o/OLiDzyFH/j6ugoqPP4mnJxqxXjXZjbUAYV8hu
3OtYr1SlNskg56+LZUdJ7k71AowbV2SEXk7zfYEqDHVDSrqNofms8BPcxG6jIlua1tWScyPkL6ui
zoNPSSvrKtNIEJNeZadGv/vczRd3zMbAy5Wm2ZMS/rJ+2JDMPHmtxZflulvcstI9wKxeP6J19jJq
vf+q6k3V7Lhw7fM0WzeOcWG51kPn6D09zc1xYTZgjXIbNBThunmGxEGDfjYIVN8C/waUxc+Z8oTK
JMY1fzXN24KOPkaKo6Fjq/vbQMHQUaeT/ALcgsJRj5p4IHTNNOuSfeKjR+ZdPh1OUCoVfOSwt0mv
Y3XyWKBa8iqCMEgVSETQ0RrNtJx+wJR9Qi3/LZRBH/vQGJ/5P1dRo4hsk9psKgwWQSMmnJMvhq2j
d7grwTFSgKhzDZ/Qk2emx+TDC9HSWNFotwvWDH9bH0G+Ik6KHQf4KkV8NcJZUyxdjRcwXu0zchAY
N6vWBME/3tqtwZyayq/PslHGvQgknI8U9aFHxqNdS42A0/7Cvqb/AKwUTU6tuo2pHsAnLt/YZ0FZ
1x3356lvdDTWQuWIRREsuVyHgNZXS69zdl4rGCUaPmLZskE1Ib6dRaZXgcTFfYRV0yMnQ/fpZpl3
M81Kh0gs5QCZGNelnzCmFSh+EBWRj13ZpKeb/xC+kZZeErqh8yOxiTThKufAb91JonuvOI3Fh7ph
5xgTIME1TfX2eDiFc4fIiPETNRBTutYSTX7xBbMhUgdMmYLAUjDuojYraxvwU97y3bhOAwRkp9q/
n4VixCWdgGrvWbZuVM5c98rvDz0GANIrtSfvVUjpx0SBYGZMrVm0im3lQmoZG5MoxToTCv+NVutm
kMw5ShJ8x8o2eVEBLb/onNeJJaBcAJYrh0OhxjunMQlpT25mSmyV+mSznrG8Me1uWaHOxE0CTh2X
SCFo9N1Gob5ksmJUkPMW77R9kT9sLSCcRiCC+pkWxQYb2aJ1vlRrAWL/oOjvch00VxFo0VCbAckg
+Idn26RT+Ruk04T/bByd7aO2gInX0aQc7VgRrP6YEjrGzwM2nPee0M0vjRPsr6dR6z6RB/7JzA2/
LTjwfyGWTPZJ4D1iKX8bjdThZ5dho0RO4ySKwKd9rTo3lh7RgVjqgveBJkbApcrLLjMJRsvY/4tU
N0yK3pBZEZIPRBCnlTR81J0AOe9U1T9hT0fHZXdCz1HQ2IMuCkk3o7oJqhhW5MZGLUzg4VBb8mo5
04xWKr03b5AZ9GpXSdY3KEfWlGDXeoyoFjaF0pcdJ6YVT8dyjlYNcr6QuuHVOEreXy7BaQZaIbXB
PtYKGXoyfUAQWQj2kCTzA/dZTnsngmjvI2ykB5ig/03F2av4P5UQc/mD5iRbgFIIUxFMH2ZVXgqB
JDmwGy+Rz4M+sNaXk1/lY0KpCmBObi49zv4vOFELiBNzYiEIPBqTPvwqWQZbDyBYB+Kq1RjoDGL4
v0bn/TiZWyJsixH1atiwkaLP/3V5FOf3fhRPpw/dWYEIj5EOWWX6IhWjB2BoZ5lLPHE5jbb+WZG4
iNvpQ7jYA+YL2JvPkAVy/tylrWTrgG2E3FQUucsY1aQvrX990WbTeDsybk2eYGGUIBJgzaYJvhtu
wgcubs5/cUDCN2Dev+9CnxSCeFwfkeke5/TzEWVjx+zFZ4z2jR/LQdmstm4V/KZQbP9IRZN/0ZSg
iJEIyxH1TKVby7UzcubUY6X+qC8kuJ7JtoZnnmUPmZ6N1paICGFVUz/N95gOq36bRjlmHlC+0dNJ
VTZYOJXxkvmF8bQt8/Q3+IVc1eAvVSaHnnE1cZICZ+mcDBH6wqXbBiD0wOy3z1I9kOPjYbxg/K7F
qlsGeLburcrmhbIj223UPH2+vPf2yV7314qv4/HaSQguCMUXfgwb1HW40m7uut4aCiFNpFBxjfQr
DExYyabZjahucHPi7zVfElmA8lyFUVMy2JFaKoNcMzI03QuMIvmeeTSfbW4WzxUVBvM2NEMKzqgm
V6lWiyWPV3qqF1e3PHCADajFSHi3lAa1DSWC9ZPHet4ODHK8dNr5AKBe5bwG8M07jco7GRJzgvQl
rYITlmSfxvFsVYCvmdaZXIkM4IbxVK1zdUv1FMxPr+WvcQ7TBKVjRj+OJvdt99DBukDzaG84mZkY
yf4Km9yPwH7zg5CIr1345Y4wTbBis1UOVvxmrt/Tr83SRiGzSYxVnyPb7mzLIVbjbWYQ/HOPPr4A
/FT8N3ImfSxg3TOdAJ7kpc0DeinDxApMWWLBTYpPfQ79rBk3oCdHdx9xzorRdnKscWARya1xdu/p
cjEn+x++etLxKFBmVQ/HcGEyr6ZHS5lNnKbuElGsgjEVJvsh0MB/o9VX0+YBCaVxvTIPPYVAtq5C
YGzxSIgTMhc8fpMqLt0Z2gqmSntniOGkx/Na1rsyufIHI5c867KAlGXHBENsZjSNTCPpINPbAKJ/
uvNVFsXf1fWixzODt17YoHj19VlnLy1Mx6V2bbOMEJiizWbg6g1H2E10qLr7u+KXQj2mkVjCa8P/
1BRhKkYuW3QQje7B7GSbUBKVoZIPXQmIRXHj+zNGriSM0NvPSJwzv4eXRLNz+yRj8wNLhRZFAyOe
VXqRJZHUfh050YdUg/NMX77s/sIKlxgihbIzV250Y92/SF9ik3TsEe3xPi82KPhrhaRTmLi2UR5k
6x8z4LrLJ4mH6MM3+8d5bezOWU5djqXCzzvsxrYsjGQNJesqx5Pies8cNM6NLBMk0pyGd8CrxFA0
6/MZ8XgHL4yjD7LtkUuvBrhmHDFWKgMqLeYYRfIWPod0hjLrQqiWLY/WtIYljVaH08HcSRyDo/aw
NhKhCNhLi0cJXX43Yvavti+gxPpXwsspk2RH0c2XieeJi61yNso2RY0UpDh+36w0JokLabI5vXwx
cSdg35f/i6S89eUMGiI9t0FWb3LO7mr6SSDsqgP8MFz6N/pbPlZsiSrwE12av67QHSRcwSpEfo1I
liXj1mygh77HA083WLttYpeyfy9n6NjtwiALfKmAaYKR0POHNlfR5VWpJs4LQd5ee0eHiFKq1z37
iSoriDTLbsFpV4Ah0rVUFi7hjzdsa0trMRF2LF3wZMvbhg+8xidQ2CSFKS/67wP/zDVi2sXBtziz
XI/P/mhxbiQXFGLTRX/k5wF3sdJA4kzJ+uHTF4hw8nqI+Zq/ofuQlGYeQY2Mg6T0pR6aAssyQjlS
AVfQYmxB3h+rK1xyRyBjzcMrniCnnnAa+FP7H9L3aqp+ETkmRCrjTnEKzaMivRl43pTTMbnbq7sk
gDenSrFSpoxCGMQtG2zyS7sx4DvNzyE3Te+LClEjqjZyrwkwKl/yYoEVcOedNYuY0tkULfAkehe4
sEVd0fasKDyWtVZ9OnSu8bTWKj+wiqWCfsDxJfiG4AQqQwXDn/ZcamoNvluodHtVO/Q0ZQMRb+jw
FW7agiEjuBFr6znk8ECNJLmLDhNJ32Yu1kpfA2YrTCdcXXLgjo0fDZirHICcgs9s6a+vNlPiim7w
AaWaOs1N7g8aNI7//fTMy7ZL+YYfJUGdxPbWYwYSGAadrzNlVWdgW4qRsfZKMkXMqYgdH/y1mRP7
xNhRtnWLhb8Uv4aImoux+xS85koziTth1nJXlm7rhQ06AYD6yxcrO/Tt3ozwS7sbAfye8yxmvvbN
SL8rA90mmJZorjIJLSno4qnc162HLYAG5Dw0HgDzMtt888kKvi05AR3yiktMQrwg1DpDwfdcgou/
QWmNOtGR3DeKnKD7vRoClrVa4SLqcuMgBWVmZRX0/tE7CIvUPZe8SJMBfKK5fIKv5/jQDcM5K+LL
`protect end_protected
